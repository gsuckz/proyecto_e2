
aaaaaaa
si