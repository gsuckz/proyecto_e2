-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Mar 21 2023 19:36:38

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top
entity top is
port (
    v_sync : out std_logic;
    pixel : out std_logic;
    led_piloto : out std_logic;
    h_sync : out std_logic;
    clk : in std_logic);
end top;

-- Architecture of top
-- View name is \INTERFACE\
architecture \INTERFACE\ of top is

signal \N__7178\ : std_logic;
signal \N__7177\ : std_logic;
signal \N__7176\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7166\ : std_logic;
signal \N__7165\ : std_logic;
signal \N__7158\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7149\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7147\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7138\ : std_logic;
signal \N__7121\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7117\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7106\ : std_logic;
signal \N__7103\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7091\ : std_logic;
signal \N__7088\ : std_logic;
signal \N__7087\ : std_logic;
signal \N__7084\ : std_logic;
signal \N__7081\ : std_logic;
signal \N__7076\ : std_logic;
signal \N__7073\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7063\ : std_logic;
signal \N__7058\ : std_logic;
signal \N__7055\ : std_logic;
signal \N__7052\ : std_logic;
signal \N__7051\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7037\ : std_logic;
signal \N__7034\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7027\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7015\ : std_logic;
signal \N__7014\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7011\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__7008\ : std_logic;
signal \N__7007\ : std_logic;
signal \N__7006\ : std_logic;
signal \N__7005\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__7002\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__7000\ : std_logic;
signal \N__6999\ : std_logic;
signal \N__6996\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6992\ : std_logic;
signal \N__6991\ : std_logic;
signal \N__6988\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6986\ : std_logic;
signal \N__6983\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6979\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6974\ : std_logic;
signal \N__6971\ : std_logic;
signal \N__6970\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6959\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6952\ : std_logic;
signal \N__6951\ : std_logic;
signal \N__6948\ : std_logic;
signal \N__6947\ : std_logic;
signal \N__6944\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6937\ : std_logic;
signal \N__6920\ : std_logic;
signal \N__6903\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6871\ : std_logic;
signal \N__6868\ : std_logic;
signal \N__6861\ : std_logic;
signal \N__6858\ : std_logic;
signal \N__6855\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6839\ : std_logic;
signal \N__6838\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6827\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6821\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6819\ : std_logic;
signal \N__6818\ : std_logic;
signal \N__6817\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6803\ : std_logic;
signal \N__6800\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6794\ : std_logic;
signal \N__6793\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6785\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6765\ : std_logic;
signal \N__6760\ : std_logic;
signal \N__6755\ : std_logic;
signal \N__6752\ : std_logic;
signal \N__6751\ : std_logic;
signal \N__6748\ : std_logic;
signal \N__6747\ : std_logic;
signal \N__6744\ : std_logic;
signal \N__6741\ : std_logic;
signal \N__6738\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6724\ : std_logic;
signal \N__6723\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6717\ : std_logic;
signal \N__6714\ : std_logic;
signal \N__6707\ : std_logic;
signal \N__6704\ : std_logic;
signal \N__6703\ : std_logic;
signal \N__6700\ : std_logic;
signal \N__6699\ : std_logic;
signal \N__6696\ : std_logic;
signal \N__6693\ : std_logic;
signal \N__6690\ : std_logic;
signal \N__6683\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6679\ : std_logic;
signal \N__6678\ : std_logic;
signal \N__6675\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6662\ : std_logic;
signal \N__6659\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6651\ : std_logic;
signal \N__6648\ : std_logic;
signal \N__6645\ : std_logic;
signal \N__6642\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6627\ : std_logic;
signal \N__6624\ : std_logic;
signal \N__6621\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6611\ : std_logic;
signal \N__6608\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6566\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6562\ : std_logic;
signal \N__6561\ : std_logic;
signal \N__6558\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6545\ : std_logic;
signal \N__6544\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6540\ : std_logic;
signal \N__6537\ : std_logic;
signal \N__6532\ : std_logic;
signal \N__6529\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6521\ : std_logic;
signal \N__6520\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6513\ : std_logic;
signal \N__6510\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6473\ : std_logic;
signal \N__6472\ : std_logic;
signal \N__6469\ : std_logic;
signal \N__6466\ : std_logic;
signal \N__6461\ : std_logic;
signal \N__6458\ : std_logic;
signal \N__6455\ : std_logic;
signal \N__6454\ : std_logic;
signal \N__6451\ : std_logic;
signal \N__6448\ : std_logic;
signal \N__6443\ : std_logic;
signal \N__6440\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6424\ : std_logic;
signal \N__6423\ : std_logic;
signal \N__6420\ : std_logic;
signal \N__6417\ : std_logic;
signal \N__6414\ : std_logic;
signal \N__6411\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6395\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6361\ : std_logic;
signal \N__6356\ : std_logic;
signal \N__6353\ : std_logic;
signal \N__6352\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6346\ : std_logic;
signal \N__6343\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6325\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6304\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6296\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6284\ : std_logic;
signal \N__6281\ : std_logic;
signal \N__6280\ : std_logic;
signal \N__6277\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6271\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6260\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6258\ : std_logic;
signal \N__6255\ : std_logic;
signal \N__6252\ : std_logic;
signal \N__6249\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6224\ : std_logic;
signal \N__6221\ : std_logic;
signal \N__6220\ : std_logic;
signal \N__6217\ : std_logic;
signal \N__6214\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6206\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6200\ : std_logic;
signal \N__6197\ : std_logic;
signal \N__6194\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6185\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6140\ : std_logic;
signal \N__6137\ : std_logic;
signal \N__6134\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6123\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__6118\ : std_logic;
signal \N__6117\ : std_logic;
signal \N__6116\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6108\ : std_logic;
signal \N__6105\ : std_logic;
signal \N__6100\ : std_logic;
signal \N__6099\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6096\ : std_logic;
signal \N__6091\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6085\ : std_logic;
signal \N__6084\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6082\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6071\ : std_logic;
signal \N__6068\ : std_logic;
signal \N__6063\ : std_logic;
signal \N__6060\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6049\ : std_logic;
signal \N__6046\ : std_logic;
signal \N__6043\ : std_logic;
signal \N__6020\ : std_logic;
signal \N__6017\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6012\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5998\ : std_logic;
signal \N__5995\ : std_logic;
signal \N__5994\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5989\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5987\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5981\ : std_logic;
signal \N__5978\ : std_logic;
signal \N__5975\ : std_logic;
signal \N__5972\ : std_logic;
signal \N__5971\ : std_logic;
signal \N__5964\ : std_logic;
signal \N__5961\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5945\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5937\ : std_logic;
signal \N__5934\ : std_logic;
signal \N__5933\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5916\ : std_logic;
signal \N__5911\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5891\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5858\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5850\ : std_logic;
signal \N__5843\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5829\ : std_logic;
signal \N__5826\ : std_logic;
signal \N__5825\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5820\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5804\ : std_logic;
signal \N__5801\ : std_logic;
signal \N__5796\ : std_logic;
signal \N__5787\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5781\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5765\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5759\ : std_logic;
signal \N__5754\ : std_logic;
signal \N__5753\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5739\ : std_logic;
signal \N__5736\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5718\ : std_logic;
signal \N__5717\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5709\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5705\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5695\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5692\ : std_logic;
signal \N__5689\ : std_logic;
signal \N__5688\ : std_logic;
signal \N__5687\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5669\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5667\ : std_logic;
signal \N__5666\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5615\ : std_logic;
signal \N__5612\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5605\ : std_logic;
signal \N__5604\ : std_logic;
signal \N__5599\ : std_logic;
signal \N__5598\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5595\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5583\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5571\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5559\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5557\ : std_logic;
signal \N__5554\ : std_logic;
signal \N__5551\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5544\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5541\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5539\ : std_logic;
signal \N__5538\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5529\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5508\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5473\ : std_logic;
signal \N__5472\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5470\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5466\ : std_logic;
signal \N__5463\ : std_logic;
signal \N__5460\ : std_logic;
signal \N__5457\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5434\ : std_logic;
signal \N__5431\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5424\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5410\ : std_logic;
signal \N__5409\ : std_logic;
signal \N__5406\ : std_logic;
signal \N__5403\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5386\ : std_logic;
signal \N__5379\ : std_logic;
signal \N__5374\ : std_logic;
signal \N__5373\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5364\ : std_logic;
signal \N__5361\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5348\ : std_logic;
signal \N__5345\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5337\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5329\ : std_logic;
signal \N__5316\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5307\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5287\ : std_logic;
signal \N__5286\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5284\ : std_logic;
signal \N__5283\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5274\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5268\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5265\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5263\ : std_logic;
signal \N__5260\ : std_logic;
signal \N__5259\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5257\ : std_logic;
signal \N__5256\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5254\ : std_logic;
signal \N__5253\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5251\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5249\ : std_logic;
signal \N__5248\ : std_logic;
signal \N__5247\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5239\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5227\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5206\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5196\ : std_logic;
signal \N__5187\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5177\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5158\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5114\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5090\ : std_logic;
signal \N__5087\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5083\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5071\ : std_logic;
signal \N__5068\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5063\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5055\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5043\ : std_logic;
signal \N__5042\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5040\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5037\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5035\ : std_logic;
signal \N__5034\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5031\ : std_logic;
signal \N__5030\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5027\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5024\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5017\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5005\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4984\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4973\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4963\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4961\ : std_logic;
signal \N__4960\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4948\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4935\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4923\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4912\ : std_logic;
signal \N__4903\ : std_logic;
signal \N__4900\ : std_logic;
signal \N__4899\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4887\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4878\ : std_logic;
signal \N__4875\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4843\ : std_logic;
signal \N__4842\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4821\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4815\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4809\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4804\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4787\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4777\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4758\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4742\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4734\ : std_logic;
signal \N__4731\ : std_logic;
signal \N__4726\ : std_logic;
signal \N__4715\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4712\ : std_logic;
signal \N__4711\ : std_logic;
signal \N__4710\ : std_logic;
signal \N__4709\ : std_logic;
signal \N__4708\ : std_logic;
signal \N__4707\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4701\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4698\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4696\ : std_logic;
signal \N__4691\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4679\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4662\ : std_logic;
signal \N__4659\ : std_logic;
signal \N__4656\ : std_logic;
signal \N__4653\ : std_logic;
signal \N__4650\ : std_logic;
signal \N__4647\ : std_logic;
signal \N__4644\ : std_logic;
signal \N__4643\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4617\ : std_logic;
signal \N__4612\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4590\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4576\ : std_logic;
signal \N__4573\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4537\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4531\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4494\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4477\ : std_logic;
signal \N__4476\ : std_logic;
signal \N__4473\ : std_logic;
signal \N__4470\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4465\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4452\ : std_logic;
signal \N__4449\ : std_logic;
signal \N__4446\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4431\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4392\ : std_logic;
signal \N__4391\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4363\ : std_logic;
signal \N__4360\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4354\ : std_logic;
signal \N__4351\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4340\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4334\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4325\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4315\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4303\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4297\ : std_logic;
signal \N__4294\ : std_logic;
signal \N__4291\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4279\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4275\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4270\ : std_logic;
signal \N__4267\ : std_logic;
signal \N__4264\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4226\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4217\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4212\ : std_logic;
signal \N__4209\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4203\ : std_logic;
signal \N__4196\ : std_logic;
signal \N__4193\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4181\ : std_logic;
signal \N__4178\ : std_logic;
signal \N__4175\ : std_logic;
signal \N__4172\ : std_logic;
signal \N__4169\ : std_logic;
signal \N__4166\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4156\ : std_logic;
signal \N__4155\ : std_logic;
signal \N__4152\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4149\ : std_logic;
signal \N__4148\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4144\ : std_logic;
signal \N__4139\ : std_logic;
signal \N__4132\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4123\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4111\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4105\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4099\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4079\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4049\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4043\ : std_logic;
signal \N__4040\ : std_logic;
signal \N__4037\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4033\ : std_logic;
signal \N__4032\ : std_logic;
signal \N__4029\ : std_logic;
signal \N__4024\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4013\ : std_logic;
signal \N__4010\ : std_logic;
signal \N__4007\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__3998\ : std_logic;
signal \N__3995\ : std_logic;
signal \N__3992\ : std_logic;
signal \N__3989\ : std_logic;
signal \N__3986\ : std_logic;
signal \N__3983\ : std_logic;
signal \N__3980\ : std_logic;
signal \N__3977\ : std_logic;
signal \N__3974\ : std_logic;
signal \N__3971\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3962\ : std_logic;
signal \N__3959\ : std_logic;
signal \N__3956\ : std_logic;
signal \N__3953\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3947\ : std_logic;
signal \N__3944\ : std_logic;
signal \N__3941\ : std_logic;
signal \N__3938\ : std_logic;
signal \N__3935\ : std_logic;
signal \N__3932\ : std_logic;
signal \N__3929\ : std_logic;
signal \N__3926\ : std_logic;
signal \N__3923\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3917\ : std_logic;
signal \N__3914\ : std_logic;
signal \N__3911\ : std_logic;
signal \N__3908\ : std_logic;
signal \N__3905\ : std_logic;
signal \N__3902\ : std_logic;
signal \N__3899\ : std_logic;
signal \N__3898\ : std_logic;
signal \N__3895\ : std_logic;
signal \N__3892\ : std_logic;
signal \N__3887\ : std_logic;
signal \N__3884\ : std_logic;
signal \N__3881\ : std_logic;
signal \N__3880\ : std_logic;
signal \N__3877\ : std_logic;
signal \N__3874\ : std_logic;
signal \N__3869\ : std_logic;
signal \N__3868\ : std_logic;
signal \N__3865\ : std_logic;
signal \N__3862\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3845\ : std_logic;
signal \N__3842\ : std_logic;
signal \N__3839\ : std_logic;
signal \N__3836\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3832\ : std_logic;
signal \N__3831\ : std_logic;
signal \N__3828\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3824\ : std_logic;
signal \N__3823\ : std_logic;
signal \N__3822\ : std_logic;
signal \N__3819\ : std_logic;
signal \N__3816\ : std_logic;
signal \N__3815\ : std_logic;
signal \N__3812\ : std_logic;
signal \N__3805\ : std_logic;
signal \N__3804\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3798\ : std_logic;
signal \N__3795\ : std_logic;
signal \N__3792\ : std_logic;
signal \N__3789\ : std_logic;
signal \N__3786\ : std_logic;
signal \N__3783\ : std_logic;
signal \N__3780\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3768\ : std_logic;
signal \N__3761\ : std_logic;
signal \N__3758\ : std_logic;
signal \N__3755\ : std_logic;
signal \N__3752\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3743\ : std_logic;
signal \N__3742\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3728\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3719\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3710\ : std_logic;
signal \N__3707\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3701\ : std_logic;
signal \N__3698\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3696\ : std_logic;
signal \N__3693\ : std_logic;
signal \N__3690\ : std_logic;
signal \N__3687\ : std_logic;
signal \N__3686\ : std_logic;
signal \N__3683\ : std_logic;
signal \N__3680\ : std_logic;
signal \N__3677\ : std_logic;
signal \N__3674\ : std_logic;
signal \N__3673\ : std_logic;
signal \N__3672\ : std_logic;
signal \N__3671\ : std_logic;
signal \N__3666\ : std_logic;
signal \N__3661\ : std_logic;
signal \N__3658\ : std_logic;
signal \N__3653\ : std_logic;
signal \N__3644\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3638\ : std_logic;
signal \N__3635\ : std_logic;
signal \N__3632\ : std_logic;
signal \N__3629\ : std_logic;
signal \N__3628\ : std_logic;
signal \N__3627\ : std_logic;
signal \N__3624\ : std_logic;
signal \N__3623\ : std_logic;
signal \N__3622\ : std_logic;
signal \N__3621\ : std_logic;
signal \N__3620\ : std_logic;
signal \N__3615\ : std_logic;
signal \N__3612\ : std_logic;
signal \N__3609\ : std_logic;
signal \N__3602\ : std_logic;
signal \N__3601\ : std_logic;
signal \N__3600\ : std_logic;
signal \N__3599\ : std_logic;
signal \N__3596\ : std_logic;
signal \N__3589\ : std_logic;
signal \N__3586\ : std_logic;
signal \N__3581\ : std_logic;
signal \N__3572\ : std_logic;
signal \N__3569\ : std_logic;
signal \N__3566\ : std_logic;
signal \N__3563\ : std_logic;
signal \N__3560\ : std_logic;
signal \N__3557\ : std_logic;
signal \N__3556\ : std_logic;
signal \N__3555\ : std_logic;
signal \N__3554\ : std_logic;
signal \N__3553\ : std_logic;
signal \N__3546\ : std_logic;
signal \N__3543\ : std_logic;
signal \N__3542\ : std_logic;
signal \N__3541\ : std_logic;
signal \N__3538\ : std_logic;
signal \N__3535\ : std_logic;
signal \N__3532\ : std_logic;
signal \N__3529\ : std_logic;
signal \N__3524\ : std_logic;
signal \N__3515\ : std_logic;
signal \N__3512\ : std_logic;
signal \N__3509\ : std_logic;
signal \N__3506\ : std_logic;
signal \N__3503\ : std_logic;
signal \N__3502\ : std_logic;
signal \N__3501\ : std_logic;
signal \N__3500\ : std_logic;
signal \N__3499\ : std_logic;
signal \N__3498\ : std_logic;
signal \N__3493\ : std_logic;
signal \N__3490\ : std_logic;
signal \N__3485\ : std_logic;
signal \N__3482\ : std_logic;
signal \N__3473\ : std_logic;
signal \N__3470\ : std_logic;
signal \N__3469\ : std_logic;
signal \N__3464\ : std_logic;
signal \N__3463\ : std_logic;
signal \N__3462\ : std_logic;
signal \N__3461\ : std_logic;
signal \N__3460\ : std_logic;
signal \N__3459\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3455\ : std_logic;
signal \N__3452\ : std_logic;
signal \N__3447\ : std_logic;
signal \N__3440\ : std_logic;
signal \N__3439\ : std_logic;
signal \N__3438\ : std_logic;
signal \N__3437\ : std_logic;
signal \N__3432\ : std_logic;
signal \N__3427\ : std_logic;
signal \N__3424\ : std_logic;
signal \N__3421\ : std_logic;
signal \N__3418\ : std_logic;
signal \N__3407\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3405\ : std_logic;
signal \N__3400\ : std_logic;
signal \N__3399\ : std_logic;
signal \N__3398\ : std_logic;
signal \N__3395\ : std_logic;
signal \N__3394\ : std_logic;
signal \N__3393\ : std_logic;
signal \N__3390\ : std_logic;
signal \N__3387\ : std_logic;
signal \N__3384\ : std_logic;
signal \N__3379\ : std_logic;
signal \N__3378\ : std_logic;
signal \N__3377\ : std_logic;
signal \N__3376\ : std_logic;
signal \N__3373\ : std_logic;
signal \N__3364\ : std_logic;
signal \N__3361\ : std_logic;
signal \N__3356\ : std_logic;
signal \N__3347\ : std_logic;
signal \N__3344\ : std_logic;
signal \N__3341\ : std_logic;
signal \N__3338\ : std_logic;
signal \N__3335\ : std_logic;
signal \N__3334\ : std_logic;
signal \N__3331\ : std_logic;
signal \N__3330\ : std_logic;
signal \N__3327\ : std_logic;
signal \N__3326\ : std_logic;
signal \N__3323\ : std_logic;
signal \N__3320\ : std_logic;
signal \N__3315\ : std_logic;
signal \N__3308\ : std_logic;
signal \N__3307\ : std_logic;
signal \N__3306\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3296\ : std_logic;
signal \N__3293\ : std_logic;
signal \N__3290\ : std_logic;
signal \N__3289\ : std_logic;
signal \N__3288\ : std_logic;
signal \N__3285\ : std_logic;
signal \N__3284\ : std_logic;
signal \N__3281\ : std_logic;
signal \N__3278\ : std_logic;
signal \N__3275\ : std_logic;
signal \N__3272\ : std_logic;
signal \N__3269\ : std_logic;
signal \N__3266\ : std_logic;
signal \N__3261\ : std_logic;
signal \N__3258\ : std_logic;
signal \N__3255\ : std_logic;
signal \N__3248\ : std_logic;
signal \N__3245\ : std_logic;
signal \N__3244\ : std_logic;
signal \N__3241\ : std_logic;
signal \N__3238\ : std_logic;
signal \N__3233\ : std_logic;
signal \N__3230\ : std_logic;
signal \N__3227\ : std_logic;
signal \N__3224\ : std_logic;
signal \N__3221\ : std_logic;
signal \N__3218\ : std_logic;
signal \N__3215\ : std_logic;
signal \N__3212\ : std_logic;
signal \N__3209\ : std_logic;
signal \N__3208\ : std_logic;
signal \N__3207\ : std_logic;
signal \N__3206\ : std_logic;
signal \N__3199\ : std_logic;
signal \N__3196\ : std_logic;
signal \N__3191\ : std_logic;
signal \N__3188\ : std_logic;
signal \N__3187\ : std_logic;
signal \N__3182\ : std_logic;
signal \N__3179\ : std_logic;
signal \N__3178\ : std_logic;
signal \N__3175\ : std_logic;
signal \N__3172\ : std_logic;
signal \N__3167\ : std_logic;
signal \N__3164\ : std_logic;
signal \N__3161\ : std_logic;
signal \N__3160\ : std_logic;
signal \N__3157\ : std_logic;
signal \N__3156\ : std_logic;
signal \N__3153\ : std_logic;
signal \N__3148\ : std_logic;
signal \N__3143\ : std_logic;
signal \N__3140\ : std_logic;
signal \N__3139\ : std_logic;
signal \N__3138\ : std_logic;
signal \N__3135\ : std_logic;
signal \N__3132\ : std_logic;
signal \N__3129\ : std_logic;
signal \N__3122\ : std_logic;
signal \N__3119\ : std_logic;
signal \N__3118\ : std_logic;
signal \N__3117\ : std_logic;
signal \N__3114\ : std_logic;
signal \N__3109\ : std_logic;
signal \N__3104\ : std_logic;
signal \N__3101\ : std_logic;
signal \N__3098\ : std_logic;
signal \N__3095\ : std_logic;
signal \N__3092\ : std_logic;
signal \N__3089\ : std_logic;
signal \N__3086\ : std_logic;
signal \N__3083\ : std_logic;
signal \N__3080\ : std_logic;
signal \N__3077\ : std_logic;
signal \N__3074\ : std_logic;
signal \N__3071\ : std_logic;
signal \N__3068\ : std_logic;
signal \N__3065\ : std_logic;
signal \N__3062\ : std_logic;
signal \N__3059\ : std_logic;
signal \N__3056\ : std_logic;
signal \N__3053\ : std_logic;
signal \N__3050\ : std_logic;
signal \N__3049\ : std_logic;
signal \N__3046\ : std_logic;
signal \N__3045\ : std_logic;
signal \N__3038\ : std_logic;
signal \N__3035\ : std_logic;
signal \N__3032\ : std_logic;
signal \N__3031\ : std_logic;
signal \N__3030\ : std_logic;
signal \N__3027\ : std_logic;
signal \N__3022\ : std_logic;
signal \N__3017\ : std_logic;
signal \N__3014\ : std_logic;
signal \N__3011\ : std_logic;
signal \N__3008\ : std_logic;
signal \N__3005\ : std_logic;
signal \N__3002\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2996\ : std_logic;
signal \N__2993\ : std_logic;
signal \N__2992\ : std_logic;
signal \N__2989\ : std_logic;
signal \N__2986\ : std_logic;
signal \N__2981\ : std_logic;
signal \N__2978\ : std_logic;
signal \N__2975\ : std_logic;
signal \N__2974\ : std_logic;
signal \N__2969\ : std_logic;
signal \N__2966\ : std_logic;
signal \N__2963\ : std_logic;
signal \N__2960\ : std_logic;
signal \N__2957\ : std_logic;
signal \N__2954\ : std_logic;
signal \N__2951\ : std_logic;
signal \N__2948\ : std_logic;
signal \N__2945\ : std_logic;
signal \N__2942\ : std_logic;
signal \N__2939\ : std_logic;
signal \N__2936\ : std_logic;
signal \N__2933\ : std_logic;
signal \N__2930\ : std_logic;
signal \N__2927\ : std_logic;
signal \N__2924\ : std_logic;
signal \N__2921\ : std_logic;
signal \N__2918\ : std_logic;
signal \N__2915\ : std_logic;
signal \N__2912\ : std_logic;
signal \N__2909\ : std_logic;
signal \N__2906\ : std_logic;
signal \N__2903\ : std_logic;
signal \N__2900\ : std_logic;
signal \N__2899\ : std_logic;
signal \N__2896\ : std_logic;
signal \N__2893\ : std_logic;
signal \N__2892\ : std_logic;
signal \N__2889\ : std_logic;
signal \N__2886\ : std_logic;
signal \N__2883\ : std_logic;
signal \N__2880\ : std_logic;
signal \N__2873\ : std_logic;
signal \N__2870\ : std_logic;
signal \N__2867\ : std_logic;
signal \N__2864\ : std_logic;
signal \N__2861\ : std_logic;
signal \N__2858\ : std_logic;
signal \N__2855\ : std_logic;
signal \N__2852\ : std_logic;
signal \N__2849\ : std_logic;
signal \N__2846\ : std_logic;
signal \N__2843\ : std_logic;
signal \N__2840\ : std_logic;
signal \N__2837\ : std_logic;
signal \N__2836\ : std_logic;
signal \N__2833\ : std_logic;
signal \N__2832\ : std_logic;
signal \N__2829\ : std_logic;
signal \N__2826\ : std_logic;
signal \N__2823\ : std_logic;
signal \N__2820\ : std_logic;
signal \N__2813\ : std_logic;
signal \N__2810\ : std_logic;
signal \N__2807\ : std_logic;
signal \N__2806\ : std_logic;
signal \N__2805\ : std_logic;
signal \N__2802\ : std_logic;
signal \N__2799\ : std_logic;
signal \N__2796\ : std_logic;
signal \N__2789\ : std_logic;
signal \N__2786\ : std_logic;
signal \N__2785\ : std_logic;
signal \N__2784\ : std_logic;
signal \N__2781\ : std_logic;
signal \N__2778\ : std_logic;
signal \N__2775\ : std_logic;
signal \N__2768\ : std_logic;
signal \N__2765\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \bfn_3_12_0_\ : std_logic;
signal \sincronismo.n1572\ : std_logic;
signal \sincronismo.n1573\ : std_logic;
signal \sincronismo.n1574\ : std_logic;
signal \sincronismo.n1575\ : std_logic;
signal \sincronismo.n1576\ : std_logic;
signal \sincronismo.n1577\ : std_logic;
signal \sincronismo.n1578\ : std_logic;
signal \sincronismo.n1579\ : std_logic;
signal \bfn_3_13_0_\ : std_logic;
signal \sincronismo.n1580\ : std_logic;
signal \sincronismo.columna_1\ : std_logic;
signal \sincronismo.columna_0\ : std_logic;
signal \sincronismo.columna_2\ : std_logic;
signal \sincronismo.n1889_cascade_\ : std_logic;
signal \sincronismo.n1193\ : std_logic;
signal h_sync_c : std_logic;
signal \sincronismo.n1383_cascade_\ : std_logic;
signal \sincronismo.n6_cascade_\ : std_logic;
signal columna_3 : std_logic;
signal n1809 : std_logic;
signal \n14_adj_131_cascade_\ : std_logic;
signal \sincronismo.n1839\ : std_logic;
signal \sincronismo.n1006_cascade_\ : std_logic;
signal \sincronismo.n10\ : std_logic;
signal \sincronismo.n1823\ : std_logic;
signal \sincronismo.n1401\ : std_logic;
signal \sincronismo.n980\ : std_logic;
signal \vsync_N_90\ : std_logic;
signal \n15_adj_136_cascade_\ : std_logic;
signal \sincronismo.n1890_cascade_\ : std_logic;
signal \sincronismo.n51\ : std_logic;
signal \salida.n1886\ : std_logic;
signal \generador.n2003_cascade_\ : std_logic;
signal \generador.px_visible_N_105_cascade_\ : std_logic;
signal pixel_c : std_logic;
signal \generador.n1856\ : std_logic;
signal \generador.n1843\ : std_logic;
signal n517 : std_logic;
signal \n1001_cascade_\ : std_logic;
signal n1167 : std_logic;
signal \generador.n6\ : std_logic;
signal linea_z_1 : std_logic;
signal \sincronismo.linea_0\ : std_logic;
signal \bfn_6_11_0_\ : std_logic;
signal \sincronismo.linea_1\ : std_logic;
signal \sincronismo.n1563\ : std_logic;
signal \sincronismo.linea_2\ : std_logic;
signal \sincronismo.n1564\ : std_logic;
signal \sincronismo.linea_3\ : std_logic;
signal \sincronismo.n1565\ : std_logic;
signal \sincronismo.n1566\ : std_logic;
signal \sincronismo.n1567\ : std_logic;
signal \sincronismo.n1568\ : std_logic;
signal \sincronismo.n1569\ : std_logic;
signal \sincronismo.n1570\ : std_logic;
signal \bfn_6_12_0_\ : std_logic;
signal \sincronismo.n1571\ : std_logic;
signal linea_9 : std_logic;
signal p_clk : std_logic;
signal \sincronismo.n1006\ : std_logic;
signal \sincronismo.n1033\ : std_logic;
signal \sincronismo.n1884\ : std_logic;
signal \sincronismo.n1932_cascade_\ : std_logic;
signal n14_adj_135 : std_logic;
signal n1928 : std_logic;
signal \n1928_cascade_\ : std_logic;
signal \n1399_cascade_\ : std_logic;
signal linea_6 : std_logic;
signal \n32_cascade_\ : std_logic;
signal \generador.n1872_cascade_\ : std_logic;
signal \generador.n1961\ : std_logic;
signal n6 : std_logic;
signal linea_7 : std_logic;
signal linea_8 : std_logic;
signal \n1946_cascade_\ : std_logic;
signal \generador.n1849\ : std_logic;
signal \n1949_cascade_\ : std_logic;
signal \generador.n1958\ : std_logic;
signal linea_5 : std_logic;
signal \generador.n2000\ : std_logic;
signal \n1363_cascade_\ : std_logic;
signal \n1955_cascade_\ : std_logic;
signal linea_4 : std_logic;
signal \generador.n1853_cascade_\ : std_logic;
signal \generador.n1855\ : std_logic;
signal \tabla.char_57_cascade_\ : std_logic;
signal \tabla.n10\ : std_logic;
signal \tabla.n10_cascade_\ : std_logic;
signal \tabla.n1365_cascade_\ : std_logic;
signal \tabla.char_6_cascade_\ : std_logic;
signal \char_code_2_cascade_\ : std_logic;
signal n1389 : std_logic;
signal n42 : std_logic;
signal \sincronismo.n1210\ : std_logic;
signal \sincronismo.n1932\ : std_logic;
signal \n1212_cascade_\ : std_logic;
signal \tabla.n7_adj_124\ : std_logic;
signal \sincronismo.n15_adj_117\ : std_logic;
signal \sincronismo.n16\ : std_logic;
signal columna_7 : std_logic;
signal \tabla.n7_adj_129\ : std_logic;
signal \tabla.n7_adj_129_cascade_\ : std_logic;
signal \tabla.char_49\ : std_logic;
signal \tabla.n7_adj_128_cascade_\ : std_logic;
signal char_42 : std_logic;
signal \generador.n1852\ : std_logic;
signal char_43 : std_logic;
signal \tabla.n728_cascade_\ : std_logic;
signal char_50 : std_logic;
signal n1952 : std_logic;
signal n58 : std_logic;
signal \n57_cascade_\ : std_logic;
signal n54 : std_logic;
signal n55 : std_logic;
signal \generador.n1964_cascade_\ : std_logic;
signal \generador.n1967\ : std_logic;
signal n1382 : std_logic;
signal \generador.n2006_cascade_\ : std_logic;
signal \generador.n1847\ : std_logic;
signal \char_13_cascade_\ : std_logic;
signal \n11_cascade_\ : std_logic;
signal \generador.n1988\ : std_logic;
signal \n1410_cascade_\ : std_logic;
signal \generador.n1991\ : std_logic;
signal \tabla.char_14_cascade_\ : std_logic;
signal n12 : std_logic;
signal \n7_cascade_\ : std_logic;
signal \n1012_cascade_\ : std_logic;
signal \generador.n1013\ : std_logic;
signal n7 : std_logic;
signal \char_5_cascade_\ : std_logic;
signal char_11 : std_logic;
signal \char_code_0_cascade_\ : std_logic;
signal \n1166_cascade_\ : std_logic;
signal \tabla.n7_adj_122_cascade_\ : std_logic;
signal \generador.n1019\ : std_logic;
signal n5 : std_logic;
signal n4 : std_logic;
signal n7_adj_137 : std_logic;
signal char_60 : std_logic;
signal n2 : std_logic;
signal \generador.n1982\ : std_logic;
signal \generador.n1985\ : std_logic;
signal \tabla.char_1\ : std_logic;
signal n1 : std_logic;
signal \generador.n1608_cascade_\ : std_logic;
signal \generador.n1008\ : std_logic;
signal \n1934_cascade_\ : std_logic;
signal \generador.n1021\ : std_logic;
signal n51 : std_logic;
signal char_61 : std_logic;
signal \tabla.n1361_cascade_\ : std_logic;
signal \n1415_cascade_\ : std_logic;
signal n1420 : std_logic;
signal \char_22_cascade_\ : std_logic;
signal \n19_cascade_\ : std_logic;
signal \tabla.n14_cascade_\ : std_logic;
signal char_20 : std_logic;
signal char_22 : std_logic;
signal n20 : std_logic;
signal n1385 : std_logic;
signal n1405 : std_logic;
signal \tabla.n7\ : std_logic;
signal n1347 : std_logic;
signal \n1347_cascade_\ : std_logic;
signal columna_8 : std_logic;
signal columna_9 : std_logic;
signal \tabla.n1930\ : std_logic;
signal \tabla.n1349\ : std_logic;
signal \tabla.n1930_cascade_\ : std_logic;
signal n1994 : std_logic;
signal \tabla.n7_adj_127\ : std_logic;
signal char_19 : std_logic;
signal columna_6 : std_logic;
signal \generador.n1976\ : std_logic;
signal \n17_cascade_\ : std_logic;
signal \generador.n1979\ : std_logic;
signal \tabla.n1397\ : std_logic;
signal n16 : std_logic;
signal n1220 : std_logic;
signal n1329 : std_logic;
signal \n1970_cascade_\ : std_logic;
signal columna_5 : std_logic;
signal \generador.n1873\ : std_logic;
signal n14_adj_133 : std_logic;
signal char_code_0 : std_logic;
signal n1166 : std_logic;
signal n1212 : std_logic;
signal \tabla.n677_cascade_\ : std_logic;
signal \tabla.char_33\ : std_logic;
signal char_code_2 : std_logic;
signal char_code_1 : std_logic;
signal n891 : std_logic;
signal char_code_3 : std_logic;
signal \tabla.n876\ : std_logic;
signal \tabla.n1361\ : std_logic;
signal \tabla.char_38\ : std_logic;
signal char_36 : std_logic;
signal char_17 : std_logic;
signal columna_4 : std_logic;
signal n24 : std_logic;
signal led_piloto_c : std_logic;
signal \n32_adj_132_cascade_\ : std_logic;
signal n31_adj_134 : std_logic;
signal n986 : std_logic;
signal \n986_cascade_\ : std_logic;
signal \n1611_cascade_\ : std_logic;
signal n38 : std_logic;
signal n33 : std_logic;
signal n35 : std_logic;
signal n34 : std_logic;
signal \n1357_cascade_\ : std_logic;
signal n1004 : std_logic;
signal \n1387_cascade_\ : std_logic;
signal \n1582_cascade_\ : std_logic;
signal n1590 : std_logic;
signal n15 : std_logic;
signal n14 : std_logic;
signal \GB_BUFFER_clk_c_THRU_CO\ : std_logic;
signal n32_adj_130 : std_logic;
signal \bfn_12_11_0_\ : std_logic;
signal n31 : std_logic;
signal n1532 : std_logic;
signal n30 : std_logic;
signal n1533 : std_logic;
signal n29 : std_logic;
signal n1534 : std_logic;
signal n28 : std_logic;
signal n1535 : std_logic;
signal n27 : std_logic;
signal n1536 : std_logic;
signal n26 : std_logic;
signal n1537 : std_logic;
signal div_led_piloto_7 : std_logic;
signal n1538 : std_logic;
signal n1539 : std_logic;
signal div_led_piloto_8 : std_logic;
signal \bfn_12_12_0_\ : std_logic;
signal div_led_piloto_9 : std_logic;
signal n1540 : std_logic;
signal div_led_piloto_10 : std_logic;
signal n1541 : std_logic;
signal div_led_piloto_11 : std_logic;
signal n1542 : std_logic;
signal div_led_piloto_12 : std_logic;
signal n1543 : std_logic;
signal div_led_piloto_13 : std_logic;
signal n1544 : std_logic;
signal div_led_piloto_14 : std_logic;
signal n1545 : std_logic;
signal div_led_piloto_15 : std_logic;
signal n1546 : std_logic;
signal n1547 : std_logic;
signal div_led_piloto_16 : std_logic;
signal \bfn_12_13_0_\ : std_logic;
signal div_led_piloto_17 : std_logic;
signal n1548 : std_logic;
signal div_led_piloto_18 : std_logic;
signal n1549 : std_logic;
signal div_led_piloto_19 : std_logic;
signal n1550 : std_logic;
signal div_led_piloto_20 : std_logic;
signal n1551 : std_logic;
signal div_led_piloto_21 : std_logic;
signal n1552 : std_logic;
signal div_led_piloto_22 : std_logic;
signal n1553 : std_logic;
signal div_led_piloto_23 : std_logic;
signal n1554 : std_logic;
signal n1555 : std_logic;
signal div_led_piloto_24 : std_logic;
signal \bfn_12_14_0_\ : std_logic;
signal div_led_piloto_25 : std_logic;
signal n1556 : std_logic;
signal div_led_piloto_26 : std_logic;
signal n1557 : std_logic;
signal div_led_piloto_27 : std_logic;
signal n1558 : std_logic;
signal div_led_piloto_28 : std_logic;
signal n1559 : std_logic;
signal div_led_piloto_29 : std_logic;
signal n1560 : std_logic;
signal div_led_piloto_30 : std_logic;
signal n1561 : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal n1562 : std_logic;
signal div_led_piloto_31 : std_logic;
signal \_gnd_net_\ : std_logic;
signal clk_c : std_logic;
signal n1029 : std_logic;

signal clk_wire : std_logic;
signal led_piloto_wire : std_logic;
signal h_sync_wire : std_logic;
signal v_sync_wire : std_logic;
signal pixel_wire : std_logic;
signal \pll.pll_px_clk_inst_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    clk_wire <= clk;
    led_piloto <= led_piloto_wire;
    h_sync <= h_sync_wire;
    v_sync <= v_sync_wire;
    pixel <= pixel_wire;
    \pll.pll_px_clk_inst_DYNAMICDELAY_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';

    \pll.pll_px_clk_inst\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "001",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0000",
            DIVQ => "101",
            DIVF => "1000010",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            LATCHINPUTVALUE => '0',
            SCLK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => OPEN,
            REFERENCECLK => \N__6401\,
            RESETB => \N__7001\,
            BYPASS => \GNDG0\,
            SDI => '0',
            DYNAMICDELAY => \pll.pll_px_clk_inst_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => p_clk
        );

    \clk_pad_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__7176\,
            GLOBALBUFFEROUTPUT => clk_c
        );

    \clk_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7178\,
            DIN => \N__7177\,
            DOUT => \N__7176\,
            PACKAGEPIN => clk_wire
        );

    \clk_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__7178\,
            PADOUT => \N__7177\,
            PADIN => \N__7176\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \led_piloto_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7167\,
            DIN => \N__7166\,
            DOUT => \N__7165\,
            PACKAGEPIN => led_piloto_wire
        );

    \led_piloto_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__7167\,
            PADOUT => \N__7166\,
            PADIN => \N__7165\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6182\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \h_sync_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7158\,
            DIN => \N__7157\,
            DOUT => \N__7156\,
            PACKAGEPIN => h_sync_wire
        );

    \h_sync_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__7158\,
            PADOUT => \N__7157\,
            PADIN => \N__7156\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2924\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \v_sync_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7149\,
            DIN => \N__7148\,
            DOUT => \N__7147\,
            PACKAGEPIN => v_sync_wire
        );

    \v_sync_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__7149\,
            PADOUT => \N__7148\,
            PADIN => \N__7147\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__2966\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \pixel_pad_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7140\,
            DIN => \N__7139\,
            DOUT => \N__7138\,
            PACKAGEPIN => pixel_wire
        );

    \pixel_pad_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__7140\,
            PADOUT => \N__7139\,
            PADIN => \N__7138\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3080\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1685\ : InMux
    port map (
            O => \N__7121\,
            I => \N__7117\
        );

    \I__1684\ : InMux
    port map (
            O => \N__7120\,
            I => \N__7114\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__7117\,
            I => div_led_piloto_25
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__7114\,
            I => div_led_piloto_25
        );

    \I__1681\ : InMux
    port map (
            O => \N__7109\,
            I => n1556
        );

    \I__1680\ : CascadeMux
    port map (
            O => \N__7106\,
            I => \N__7103\
        );

    \I__1679\ : InMux
    port map (
            O => \N__7103\,
            I => \N__7099\
        );

    \I__1678\ : InMux
    port map (
            O => \N__7102\,
            I => \N__7096\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__7099\,
            I => div_led_piloto_26
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__7096\,
            I => div_led_piloto_26
        );

    \I__1675\ : InMux
    port map (
            O => \N__7091\,
            I => n1557
        );

    \I__1674\ : InMux
    port map (
            O => \N__7088\,
            I => \N__7084\
        );

    \I__1673\ : InMux
    port map (
            O => \N__7087\,
            I => \N__7081\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__7084\,
            I => div_led_piloto_27
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__7081\,
            I => div_led_piloto_27
        );

    \I__1670\ : InMux
    port map (
            O => \N__7076\,
            I => n1558
        );

    \I__1669\ : CascadeMux
    port map (
            O => \N__7073\,
            I => \N__7070\
        );

    \I__1668\ : InMux
    port map (
            O => \N__7070\,
            I => \N__7066\
        );

    \I__1667\ : InMux
    port map (
            O => \N__7069\,
            I => \N__7063\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__7066\,
            I => div_led_piloto_28
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__7063\,
            I => div_led_piloto_28
        );

    \I__1664\ : InMux
    port map (
            O => \N__7058\,
            I => n1559
        );

    \I__1663\ : InMux
    port map (
            O => \N__7055\,
            I => \N__7052\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__7052\,
            I => \N__7048\
        );

    \I__1661\ : InMux
    port map (
            O => \N__7051\,
            I => \N__7045\
        );

    \I__1660\ : Span4Mux_h
    port map (
            O => \N__7048\,
            I => \N__7042\
        );

    \I__1659\ : LocalMux
    port map (
            O => \N__7045\,
            I => div_led_piloto_29
        );

    \I__1658\ : Odrv4
    port map (
            O => \N__7042\,
            I => div_led_piloto_29
        );

    \I__1657\ : InMux
    port map (
            O => \N__7037\,
            I => n1560
        );

    \I__1656\ : CascadeMux
    port map (
            O => \N__7034\,
            I => \N__7031\
        );

    \I__1655\ : InMux
    port map (
            O => \N__7031\,
            I => \N__7027\
        );

    \I__1654\ : InMux
    port map (
            O => \N__7030\,
            I => \N__7024\
        );

    \I__1653\ : LocalMux
    port map (
            O => \N__7027\,
            I => div_led_piloto_30
        );

    \I__1652\ : LocalMux
    port map (
            O => \N__7024\,
            I => div_led_piloto_30
        );

    \I__1651\ : InMux
    port map (
            O => \N__7019\,
            I => n1561
        );

    \I__1650\ : CascadeMux
    port map (
            O => \N__7016\,
            I => \N__6996\
        );

    \I__1649\ : CascadeMux
    port map (
            O => \N__7015\,
            I => \N__6992\
        );

    \I__1648\ : CascadeMux
    port map (
            O => \N__7014\,
            I => \N__6988\
        );

    \I__1647\ : CascadeMux
    port map (
            O => \N__7013\,
            I => \N__6983\
        );

    \I__1646\ : CascadeMux
    port map (
            O => \N__7012\,
            I => \N__6979\
        );

    \I__1645\ : CascadeMux
    port map (
            O => \N__7011\,
            I => \N__6975\
        );

    \I__1644\ : CascadeMux
    port map (
            O => \N__7010\,
            I => \N__6971\
        );

    \I__1643\ : CascadeMux
    port map (
            O => \N__7009\,
            I => \N__6967\
        );

    \I__1642\ : CascadeMux
    port map (
            O => \N__7008\,
            I => \N__6963\
        );

    \I__1641\ : CascadeMux
    port map (
            O => \N__7007\,
            I => \N__6959\
        );

    \I__1640\ : CascadeMux
    port map (
            O => \N__7006\,
            I => \N__6955\
        );

    \I__1639\ : CascadeMux
    port map (
            O => \N__7005\,
            I => \N__6952\
        );

    \I__1638\ : CascadeMux
    port map (
            O => \N__7004\,
            I => \N__6948\
        );

    \I__1637\ : CascadeMux
    port map (
            O => \N__7003\,
            I => \N__6944\
        );

    \I__1636\ : CascadeMux
    port map (
            O => \N__7002\,
            I => \N__6940\
        );

    \I__1635\ : IoInMux
    port map (
            O => \N__7001\,
            I => \N__6937\
        );

    \I__1634\ : InMux
    port map (
            O => \N__7000\,
            I => \N__6920\
        );

    \I__1633\ : InMux
    port map (
            O => \N__6999\,
            I => \N__6920\
        );

    \I__1632\ : InMux
    port map (
            O => \N__6996\,
            I => \N__6920\
        );

    \I__1631\ : InMux
    port map (
            O => \N__6995\,
            I => \N__6920\
        );

    \I__1630\ : InMux
    port map (
            O => \N__6992\,
            I => \N__6920\
        );

    \I__1629\ : InMux
    port map (
            O => \N__6991\,
            I => \N__6920\
        );

    \I__1628\ : InMux
    port map (
            O => \N__6988\,
            I => \N__6920\
        );

    \I__1627\ : InMux
    port map (
            O => \N__6987\,
            I => \N__6920\
        );

    \I__1626\ : InMux
    port map (
            O => \N__6986\,
            I => \N__6903\
        );

    \I__1625\ : InMux
    port map (
            O => \N__6983\,
            I => \N__6903\
        );

    \I__1624\ : InMux
    port map (
            O => \N__6982\,
            I => \N__6903\
        );

    \I__1623\ : InMux
    port map (
            O => \N__6979\,
            I => \N__6903\
        );

    \I__1622\ : InMux
    port map (
            O => \N__6978\,
            I => \N__6903\
        );

    \I__1621\ : InMux
    port map (
            O => \N__6975\,
            I => \N__6903\
        );

    \I__1620\ : InMux
    port map (
            O => \N__6974\,
            I => \N__6903\
        );

    \I__1619\ : InMux
    port map (
            O => \N__6971\,
            I => \N__6903\
        );

    \I__1618\ : InMux
    port map (
            O => \N__6970\,
            I => \N__6886\
        );

    \I__1617\ : InMux
    port map (
            O => \N__6967\,
            I => \N__6886\
        );

    \I__1616\ : InMux
    port map (
            O => \N__6966\,
            I => \N__6886\
        );

    \I__1615\ : InMux
    port map (
            O => \N__6963\,
            I => \N__6886\
        );

    \I__1614\ : InMux
    port map (
            O => \N__6962\,
            I => \N__6886\
        );

    \I__1613\ : InMux
    port map (
            O => \N__6959\,
            I => \N__6886\
        );

    \I__1612\ : InMux
    port map (
            O => \N__6958\,
            I => \N__6886\
        );

    \I__1611\ : InMux
    port map (
            O => \N__6955\,
            I => \N__6886\
        );

    \I__1610\ : InMux
    port map (
            O => \N__6952\,
            I => \N__6871\
        );

    \I__1609\ : InMux
    port map (
            O => \N__6951\,
            I => \N__6871\
        );

    \I__1608\ : InMux
    port map (
            O => \N__6948\,
            I => \N__6871\
        );

    \I__1607\ : InMux
    port map (
            O => \N__6947\,
            I => \N__6871\
        );

    \I__1606\ : InMux
    port map (
            O => \N__6944\,
            I => \N__6871\
        );

    \I__1605\ : InMux
    port map (
            O => \N__6943\,
            I => \N__6871\
        );

    \I__1604\ : InMux
    port map (
            O => \N__6940\,
            I => \N__6871\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__6937\,
            I => \N__6868\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__6920\,
            I => \N__6861\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__6903\,
            I => \N__6861\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__6886\,
            I => \N__6861\
        );

    \I__1599\ : LocalMux
    port map (
            O => \N__6871\,
            I => \N__6858\
        );

    \I__1598\ : Span4Mux_s2_v
    port map (
            O => \N__6868\,
            I => \N__6855\
        );

    \I__1597\ : Span12Mux_v
    port map (
            O => \N__6861\,
            I => \N__6850\
        );

    \I__1596\ : Sp12to4
    port map (
            O => \N__6858\,
            I => \N__6850\
        );

    \I__1595\ : Span4Mux_v
    port map (
            O => \N__6855\,
            I => \N__6847\
        );

    \I__1594\ : Odrv12
    port map (
            O => \N__6850\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1593\ : Odrv4
    port map (
            O => \N__6847\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1592\ : InMux
    port map (
            O => \N__6842\,
            I => n1562
        );

    \I__1591\ : InMux
    port map (
            O => \N__6839\,
            I => \N__6835\
        );

    \I__1590\ : InMux
    port map (
            O => \N__6838\,
            I => \N__6832\
        );

    \I__1589\ : LocalMux
    port map (
            O => \N__6835\,
            I => div_led_piloto_31
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__6832\,
            I => div_led_piloto_31
        );

    \I__1587\ : InMux
    port map (
            O => \N__6827\,
            I => \N__6824\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__6824\,
            I => \N__6821\
        );

    \I__1585\ : Glb2LocalMux
    port map (
            O => \N__6821\,
            I => \N__6806\
        );

    \I__1584\ : ClkMux
    port map (
            O => \N__6820\,
            I => \N__6806\
        );

    \I__1583\ : ClkMux
    port map (
            O => \N__6819\,
            I => \N__6806\
        );

    \I__1582\ : ClkMux
    port map (
            O => \N__6818\,
            I => \N__6806\
        );

    \I__1581\ : ClkMux
    port map (
            O => \N__6817\,
            I => \N__6806\
        );

    \I__1580\ : GlobalMux
    port map (
            O => \N__6806\,
            I => \N__6803\
        );

    \I__1579\ : gio2CtrlBuf
    port map (
            O => \N__6803\,
            I => clk_c
        );

    \I__1578\ : SRMux
    port map (
            O => \N__6800\,
            I => \N__6797\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__6797\,
            I => \N__6794\
        );

    \I__1576\ : Span4Mux_h
    port map (
            O => \N__6794\,
            I => \N__6788\
        );

    \I__1575\ : SRMux
    port map (
            O => \N__6793\,
            I => \N__6785\
        );

    \I__1574\ : SRMux
    port map (
            O => \N__6792\,
            I => \N__6782\
        );

    \I__1573\ : SRMux
    port map (
            O => \N__6791\,
            I => \N__6779\
        );

    \I__1572\ : Odrv4
    port map (
            O => \N__6788\,
            I => n1029
        );

    \I__1571\ : LocalMux
    port map (
            O => \N__6785\,
            I => n1029
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__6782\,
            I => n1029
        );

    \I__1569\ : LocalMux
    port map (
            O => \N__6779\,
            I => n1029
        );

    \I__1568\ : InMux
    port map (
            O => \N__6770\,
            I => \N__6765\
        );

    \I__1567\ : InMux
    port map (
            O => \N__6769\,
            I => \N__6760\
        );

    \I__1566\ : InMux
    port map (
            O => \N__6768\,
            I => \N__6760\
        );

    \I__1565\ : LocalMux
    port map (
            O => \N__6765\,
            I => div_led_piloto_16
        );

    \I__1564\ : LocalMux
    port map (
            O => \N__6760\,
            I => div_led_piloto_16
        );

    \I__1563\ : InMux
    port map (
            O => \N__6755\,
            I => \bfn_12_13_0_\
        );

    \I__1562\ : CascadeMux
    port map (
            O => \N__6752\,
            I => \N__6748\
        );

    \I__1561\ : InMux
    port map (
            O => \N__6751\,
            I => \N__6744\
        );

    \I__1560\ : InMux
    port map (
            O => \N__6748\,
            I => \N__6741\
        );

    \I__1559\ : InMux
    port map (
            O => \N__6747\,
            I => \N__6738\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__6744\,
            I => div_led_piloto_17
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__6741\,
            I => div_led_piloto_17
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__6738\,
            I => div_led_piloto_17
        );

    \I__1555\ : InMux
    port map (
            O => \N__6731\,
            I => n1548
        );

    \I__1554\ : InMux
    port map (
            O => \N__6728\,
            I => \N__6725\
        );

    \I__1553\ : LocalMux
    port map (
            O => \N__6725\,
            I => \N__6720\
        );

    \I__1552\ : InMux
    port map (
            O => \N__6724\,
            I => \N__6717\
        );

    \I__1551\ : InMux
    port map (
            O => \N__6723\,
            I => \N__6714\
        );

    \I__1550\ : Odrv4
    port map (
            O => \N__6720\,
            I => div_led_piloto_18
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__6717\,
            I => div_led_piloto_18
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__6714\,
            I => div_led_piloto_18
        );

    \I__1547\ : InMux
    port map (
            O => \N__6707\,
            I => n1549
        );

    \I__1546\ : CascadeMux
    port map (
            O => \N__6704\,
            I => \N__6700\
        );

    \I__1545\ : InMux
    port map (
            O => \N__6703\,
            I => \N__6696\
        );

    \I__1544\ : InMux
    port map (
            O => \N__6700\,
            I => \N__6693\
        );

    \I__1543\ : InMux
    port map (
            O => \N__6699\,
            I => \N__6690\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__6696\,
            I => div_led_piloto_19
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__6693\,
            I => div_led_piloto_19
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__6690\,
            I => div_led_piloto_19
        );

    \I__1539\ : InMux
    port map (
            O => \N__6683\,
            I => n1550
        );

    \I__1538\ : InMux
    port map (
            O => \N__6680\,
            I => \N__6675\
        );

    \I__1537\ : InMux
    port map (
            O => \N__6679\,
            I => \N__6672\
        );

    \I__1536\ : InMux
    port map (
            O => \N__6678\,
            I => \N__6669\
        );

    \I__1535\ : LocalMux
    port map (
            O => \N__6675\,
            I => div_led_piloto_20
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__6672\,
            I => div_led_piloto_20
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__6669\,
            I => div_led_piloto_20
        );

    \I__1532\ : InMux
    port map (
            O => \N__6662\,
            I => n1551
        );

    \I__1531\ : InMux
    port map (
            O => \N__6659\,
            I => \N__6655\
        );

    \I__1530\ : CascadeMux
    port map (
            O => \N__6658\,
            I => \N__6652\
        );

    \I__1529\ : LocalMux
    port map (
            O => \N__6655\,
            I => \N__6648\
        );

    \I__1528\ : InMux
    port map (
            O => \N__6652\,
            I => \N__6645\
        );

    \I__1527\ : InMux
    port map (
            O => \N__6651\,
            I => \N__6642\
        );

    \I__1526\ : Odrv4
    port map (
            O => \N__6648\,
            I => div_led_piloto_21
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__6645\,
            I => div_led_piloto_21
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__6642\,
            I => div_led_piloto_21
        );

    \I__1523\ : InMux
    port map (
            O => \N__6635\,
            I => n1552
        );

    \I__1522\ : InMux
    port map (
            O => \N__6632\,
            I => \N__6629\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__6629\,
            I => \N__6624\
        );

    \I__1520\ : InMux
    port map (
            O => \N__6628\,
            I => \N__6621\
        );

    \I__1519\ : InMux
    port map (
            O => \N__6627\,
            I => \N__6618\
        );

    \I__1518\ : Odrv4
    port map (
            O => \N__6624\,
            I => div_led_piloto_22
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__6621\,
            I => div_led_piloto_22
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__6618\,
            I => div_led_piloto_22
        );

    \I__1515\ : InMux
    port map (
            O => \N__6611\,
            I => n1553
        );

    \I__1514\ : CascadeMux
    port map (
            O => \N__6608\,
            I => \N__6604\
        );

    \I__1513\ : CascadeMux
    port map (
            O => \N__6607\,
            I => \N__6601\
        );

    \I__1512\ : InMux
    port map (
            O => \N__6604\,
            I => \N__6598\
        );

    \I__1511\ : InMux
    port map (
            O => \N__6601\,
            I => \N__6595\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__6598\,
            I => div_led_piloto_23
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__6595\,
            I => div_led_piloto_23
        );

    \I__1508\ : InMux
    port map (
            O => \N__6590\,
            I => n1554
        );

    \I__1507\ : CascadeMux
    port map (
            O => \N__6587\,
            I => \N__6583\
        );

    \I__1506\ : CascadeMux
    port map (
            O => \N__6586\,
            I => \N__6580\
        );

    \I__1505\ : InMux
    port map (
            O => \N__6583\,
            I => \N__6577\
        );

    \I__1504\ : InMux
    port map (
            O => \N__6580\,
            I => \N__6574\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__6577\,
            I => \N__6571\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__6574\,
            I => div_led_piloto_24
        );

    \I__1501\ : Odrv4
    port map (
            O => \N__6571\,
            I => div_led_piloto_24
        );

    \I__1500\ : InMux
    port map (
            O => \N__6566\,
            I => \bfn_12_14_0_\
        );

    \I__1499\ : InMux
    port map (
            O => \N__6563\,
            I => \N__6558\
        );

    \I__1498\ : InMux
    port map (
            O => \N__6562\,
            I => \N__6553\
        );

    \I__1497\ : InMux
    port map (
            O => \N__6561\,
            I => \N__6553\
        );

    \I__1496\ : LocalMux
    port map (
            O => \N__6558\,
            I => div_led_piloto_8
        );

    \I__1495\ : LocalMux
    port map (
            O => \N__6553\,
            I => div_led_piloto_8
        );

    \I__1494\ : InMux
    port map (
            O => \N__6548\,
            I => \bfn_12_12_0_\
        );

    \I__1493\ : CascadeMux
    port map (
            O => \N__6545\,
            I => \N__6540\
        );

    \I__1492\ : CascadeMux
    port map (
            O => \N__6544\,
            I => \N__6537\
        );

    \I__1491\ : InMux
    port map (
            O => \N__6543\,
            I => \N__6532\
        );

    \I__1490\ : InMux
    port map (
            O => \N__6540\,
            I => \N__6532\
        );

    \I__1489\ : InMux
    port map (
            O => \N__6537\,
            I => \N__6529\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__6532\,
            I => div_led_piloto_9
        );

    \I__1487\ : LocalMux
    port map (
            O => \N__6529\,
            I => div_led_piloto_9
        );

    \I__1486\ : InMux
    port map (
            O => \N__6524\,
            I => n1540
        );

    \I__1485\ : InMux
    port map (
            O => \N__6521\,
            I => \N__6516\
        );

    \I__1484\ : InMux
    port map (
            O => \N__6520\,
            I => \N__6513\
        );

    \I__1483\ : InMux
    port map (
            O => \N__6519\,
            I => \N__6510\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__6516\,
            I => div_led_piloto_10
        );

    \I__1481\ : LocalMux
    port map (
            O => \N__6513\,
            I => div_led_piloto_10
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__6510\,
            I => div_led_piloto_10
        );

    \I__1479\ : InMux
    port map (
            O => \N__6503\,
            I => n1541
        );

    \I__1478\ : CascadeMux
    port map (
            O => \N__6500\,
            I => \N__6495\
        );

    \I__1477\ : CascadeMux
    port map (
            O => \N__6499\,
            I => \N__6492\
        );

    \I__1476\ : InMux
    port map (
            O => \N__6498\,
            I => \N__6489\
        );

    \I__1475\ : InMux
    port map (
            O => \N__6495\,
            I => \N__6486\
        );

    \I__1474\ : InMux
    port map (
            O => \N__6492\,
            I => \N__6483\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__6489\,
            I => div_led_piloto_11
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__6486\,
            I => div_led_piloto_11
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__6483\,
            I => div_led_piloto_11
        );

    \I__1470\ : InMux
    port map (
            O => \N__6476\,
            I => n1542
        );

    \I__1469\ : InMux
    port map (
            O => \N__6473\,
            I => \N__6469\
        );

    \I__1468\ : InMux
    port map (
            O => \N__6472\,
            I => \N__6466\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__6469\,
            I => div_led_piloto_12
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__6466\,
            I => div_led_piloto_12
        );

    \I__1465\ : InMux
    port map (
            O => \N__6461\,
            I => n1543
        );

    \I__1464\ : CascadeMux
    port map (
            O => \N__6458\,
            I => \N__6455\
        );

    \I__1463\ : InMux
    port map (
            O => \N__6455\,
            I => \N__6451\
        );

    \I__1462\ : InMux
    port map (
            O => \N__6454\,
            I => \N__6448\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__6451\,
            I => div_led_piloto_13
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__6448\,
            I => div_led_piloto_13
        );

    \I__1459\ : InMux
    port map (
            O => \N__6443\,
            I => n1544
        );

    \I__1458\ : InMux
    port map (
            O => \N__6440\,
            I => \N__6436\
        );

    \I__1457\ : InMux
    port map (
            O => \N__6439\,
            I => \N__6433\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__6436\,
            I => div_led_piloto_14
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__6433\,
            I => div_led_piloto_14
        );

    \I__1454\ : InMux
    port map (
            O => \N__6428\,
            I => n1545
        );

    \I__1453\ : CascadeMux
    port map (
            O => \N__6425\,
            I => \N__6420\
        );

    \I__1452\ : InMux
    port map (
            O => \N__6424\,
            I => \N__6417\
        );

    \I__1451\ : InMux
    port map (
            O => \N__6423\,
            I => \N__6414\
        );

    \I__1450\ : InMux
    port map (
            O => \N__6420\,
            I => \N__6411\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__6417\,
            I => div_led_piloto_15
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__6414\,
            I => div_led_piloto_15
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__6411\,
            I => div_led_piloto_15
        );

    \I__1446\ : InMux
    port map (
            O => \N__6404\,
            I => n1546
        );

    \I__1445\ : IoInMux
    port map (
            O => \N__6401\,
            I => \N__6398\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__6398\,
            I => \N__6395\
        );

    \I__1443\ : Span4Mux_s2_v
    port map (
            O => \N__6395\,
            I => \N__6392\
        );

    \I__1442\ : Span4Mux_v
    port map (
            O => \N__6392\,
            I => \N__6389\
        );

    \I__1441\ : Odrv4
    port map (
            O => \N__6389\,
            I => \GB_BUFFER_clk_c_THRU_CO\
        );

    \I__1440\ : InMux
    port map (
            O => \N__6386\,
            I => \N__6382\
        );

    \I__1439\ : InMux
    port map (
            O => \N__6385\,
            I => \N__6379\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__6382\,
            I => n32_adj_130
        );

    \I__1437\ : LocalMux
    port map (
            O => \N__6379\,
            I => n32_adj_130
        );

    \I__1436\ : InMux
    port map (
            O => \N__6374\,
            I => \bfn_12_11_0_\
        );

    \I__1435\ : CascadeMux
    port map (
            O => \N__6371\,
            I => \N__6367\
        );

    \I__1434\ : InMux
    port map (
            O => \N__6370\,
            I => \N__6364\
        );

    \I__1433\ : InMux
    port map (
            O => \N__6367\,
            I => \N__6361\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__6364\,
            I => n31
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__6361\,
            I => n31
        );

    \I__1430\ : InMux
    port map (
            O => \N__6356\,
            I => n1532
        );

    \I__1429\ : CascadeMux
    port map (
            O => \N__6353\,
            I => \N__6349\
        );

    \I__1428\ : InMux
    port map (
            O => \N__6352\,
            I => \N__6346\
        );

    \I__1427\ : InMux
    port map (
            O => \N__6349\,
            I => \N__6343\
        );

    \I__1426\ : LocalMux
    port map (
            O => \N__6346\,
            I => n30
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__6343\,
            I => n30
        );

    \I__1424\ : InMux
    port map (
            O => \N__6338\,
            I => n1533
        );

    \I__1423\ : CascadeMux
    port map (
            O => \N__6335\,
            I => \N__6331\
        );

    \I__1422\ : InMux
    port map (
            O => \N__6334\,
            I => \N__6328\
        );

    \I__1421\ : InMux
    port map (
            O => \N__6331\,
            I => \N__6325\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__6328\,
            I => n29
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__6325\,
            I => n29
        );

    \I__1418\ : InMux
    port map (
            O => \N__6320\,
            I => n1534
        );

    \I__1417\ : CascadeMux
    port map (
            O => \N__6317\,
            I => \N__6313\
        );

    \I__1416\ : CascadeMux
    port map (
            O => \N__6316\,
            I => \N__6310\
        );

    \I__1415\ : InMux
    port map (
            O => \N__6313\,
            I => \N__6307\
        );

    \I__1414\ : InMux
    port map (
            O => \N__6310\,
            I => \N__6304\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__6307\,
            I => n28
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__6304\,
            I => n28
        );

    \I__1411\ : InMux
    port map (
            O => \N__6299\,
            I => n1535
        );

    \I__1410\ : InMux
    port map (
            O => \N__6296\,
            I => \N__6292\
        );

    \I__1409\ : InMux
    port map (
            O => \N__6295\,
            I => \N__6289\
        );

    \I__1408\ : LocalMux
    port map (
            O => \N__6292\,
            I => n27
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__6289\,
            I => n27
        );

    \I__1406\ : InMux
    port map (
            O => \N__6284\,
            I => n1536
        );

    \I__1405\ : CascadeMux
    port map (
            O => \N__6281\,
            I => \N__6277\
        );

    \I__1404\ : InMux
    port map (
            O => \N__6280\,
            I => \N__6274\
        );

    \I__1403\ : InMux
    port map (
            O => \N__6277\,
            I => \N__6271\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__6274\,
            I => n26
        );

    \I__1401\ : LocalMux
    port map (
            O => \N__6271\,
            I => n26
        );

    \I__1400\ : InMux
    port map (
            O => \N__6266\,
            I => n1537
        );

    \I__1399\ : InMux
    port map (
            O => \N__6263\,
            I => \N__6260\
        );

    \I__1398\ : LocalMux
    port map (
            O => \N__6260\,
            I => \N__6255\
        );

    \I__1397\ : InMux
    port map (
            O => \N__6259\,
            I => \N__6252\
        );

    \I__1396\ : InMux
    port map (
            O => \N__6258\,
            I => \N__6249\
        );

    \I__1395\ : Odrv4
    port map (
            O => \N__6255\,
            I => div_led_piloto_7
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__6252\,
            I => div_led_piloto_7
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__6249\,
            I => div_led_piloto_7
        );

    \I__1392\ : InMux
    port map (
            O => \N__6242\,
            I => n1538
        );

    \I__1391\ : InMux
    port map (
            O => \N__6239\,
            I => \N__6236\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__6236\,
            I => n35
        );

    \I__1389\ : InMux
    port map (
            O => \N__6233\,
            I => \N__6230\
        );

    \I__1388\ : LocalMux
    port map (
            O => \N__6230\,
            I => n34
        );

    \I__1387\ : CascadeMux
    port map (
            O => \N__6227\,
            I => \n1357_cascade_\
        );

    \I__1386\ : InMux
    port map (
            O => \N__6224\,
            I => \N__6221\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__6221\,
            I => \N__6217\
        );

    \I__1384\ : InMux
    port map (
            O => \N__6220\,
            I => \N__6214\
        );

    \I__1383\ : Odrv4
    port map (
            O => \N__6217\,
            I => n1004
        );

    \I__1382\ : LocalMux
    port map (
            O => \N__6214\,
            I => n1004
        );

    \I__1381\ : CascadeMux
    port map (
            O => \N__6209\,
            I => \n1387_cascade_\
        );

    \I__1380\ : CascadeMux
    port map (
            O => \N__6206\,
            I => \n1582_cascade_\
        );

    \I__1379\ : CascadeMux
    port map (
            O => \N__6203\,
            I => \N__6200\
        );

    \I__1378\ : InMux
    port map (
            O => \N__6200\,
            I => \N__6197\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__6197\,
            I => n1590
        );

    \I__1376\ : InMux
    port map (
            O => \N__6194\,
            I => \N__6191\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__6191\,
            I => n15
        );

    \I__1374\ : InMux
    port map (
            O => \N__6188\,
            I => \N__6185\
        );

    \I__1373\ : LocalMux
    port map (
            O => \N__6185\,
            I => n14
        );

    \I__1372\ : IoInMux
    port map (
            O => \N__6182\,
            I => \N__6179\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__6179\,
            I => \N__6176\
        );

    \I__1370\ : Span4Mux_s0_h
    port map (
            O => \N__6176\,
            I => \N__6173\
        );

    \I__1369\ : Sp12to4
    port map (
            O => \N__6173\,
            I => \N__6170\
        );

    \I__1368\ : Span12Mux_v
    port map (
            O => \N__6170\,
            I => \N__6167\
        );

    \I__1367\ : Span12Mux_h
    port map (
            O => \N__6167\,
            I => \N__6164\
        );

    \I__1366\ : Odrv12
    port map (
            O => \N__6164\,
            I => led_piloto_c
        );

    \I__1365\ : CascadeMux
    port map (
            O => \N__6161\,
            I => \n32_adj_132_cascade_\
        );

    \I__1364\ : InMux
    port map (
            O => \N__6158\,
            I => \N__6155\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__6155\,
            I => n31_adj_134
        );

    \I__1362\ : InMux
    port map (
            O => \N__6152\,
            I => \N__6149\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__6149\,
            I => n986
        );

    \I__1360\ : CascadeMux
    port map (
            O => \N__6146\,
            I => \n986_cascade_\
        );

    \I__1359\ : CascadeMux
    port map (
            O => \N__6143\,
            I => \n1611_cascade_\
        );

    \I__1358\ : InMux
    port map (
            O => \N__6140\,
            I => \N__6137\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__6137\,
            I => n38
        );

    \I__1356\ : InMux
    port map (
            O => \N__6134\,
            I => \N__6131\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__6131\,
            I => n33
        );

    \I__1354\ : InMux
    port map (
            O => \N__6128\,
            I => \N__6124\
        );

    \I__1353\ : InMux
    port map (
            O => \N__6127\,
            I => \N__6120\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__6124\,
            I => \N__6111\
        );

    \I__1351\ : InMux
    port map (
            O => \N__6123\,
            I => \N__6108\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__6120\,
            I => \N__6105\
        );

    \I__1349\ : InMux
    port map (
            O => \N__6119\,
            I => \N__6100\
        );

    \I__1348\ : InMux
    port map (
            O => \N__6118\,
            I => \N__6100\
        );

    \I__1347\ : InMux
    port map (
            O => \N__6117\,
            I => \N__6091\
        );

    \I__1346\ : InMux
    port map (
            O => \N__6116\,
            I => \N__6091\
        );

    \I__1345\ : InMux
    port map (
            O => \N__6115\,
            I => \N__6088\
        );

    \I__1344\ : InMux
    port map (
            O => \N__6114\,
            I => \N__6085\
        );

    \I__1343\ : Span4Mux_v
    port map (
            O => \N__6111\,
            I => \N__6079\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__6108\,
            I => \N__6076\
        );

    \I__1341\ : Span4Mux_h
    port map (
            O => \N__6105\,
            I => \N__6071\
        );

    \I__1340\ : LocalMux
    port map (
            O => \N__6100\,
            I => \N__6071\
        );

    \I__1339\ : InMux
    port map (
            O => \N__6099\,
            I => \N__6068\
        );

    \I__1338\ : InMux
    port map (
            O => \N__6098\,
            I => \N__6063\
        );

    \I__1337\ : InMux
    port map (
            O => \N__6097\,
            I => \N__6063\
        );

    \I__1336\ : InMux
    port map (
            O => \N__6096\,
            I => \N__6060\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__6091\,
            I => \N__6055\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__6088\,
            I => \N__6055\
        );

    \I__1333\ : LocalMux
    port map (
            O => \N__6085\,
            I => \N__6052\
        );

    \I__1332\ : InMux
    port map (
            O => \N__6084\,
            I => \N__6049\
        );

    \I__1331\ : InMux
    port map (
            O => \N__6083\,
            I => \N__6046\
        );

    \I__1330\ : InMux
    port map (
            O => \N__6082\,
            I => \N__6043\
        );

    \I__1329\ : Odrv4
    port map (
            O => \N__6079\,
            I => n1329
        );

    \I__1328\ : Odrv4
    port map (
            O => \N__6076\,
            I => n1329
        );

    \I__1327\ : Odrv4
    port map (
            O => \N__6071\,
            I => n1329
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__6068\,
            I => n1329
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__6063\,
            I => n1329
        );

    \I__1324\ : LocalMux
    port map (
            O => \N__6060\,
            I => n1329
        );

    \I__1323\ : Odrv4
    port map (
            O => \N__6055\,
            I => n1329
        );

    \I__1322\ : Odrv12
    port map (
            O => \N__6052\,
            I => n1329
        );

    \I__1321\ : LocalMux
    port map (
            O => \N__6049\,
            I => n1329
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__6046\,
            I => n1329
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__6043\,
            I => n1329
        );

    \I__1318\ : CascadeMux
    port map (
            O => \N__6020\,
            I => \n1970_cascade_\
        );

    \I__1317\ : InMux
    port map (
            O => \N__6017\,
            I => \N__6007\
        );

    \I__1316\ : InMux
    port map (
            O => \N__6016\,
            I => \N__6007\
        );

    \I__1315\ : InMux
    port map (
            O => \N__6015\,
            I => \N__6004\
        );

    \I__1314\ : InMux
    port map (
            O => \N__6014\,
            I => \N__6001\
        );

    \I__1313\ : InMux
    port map (
            O => \N__6013\,
            I => \N__5998\
        );

    \I__1312\ : CascadeMux
    port map (
            O => \N__6012\,
            I => \N__5995\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__6007\,
            I => \N__5984\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__6004\,
            I => \N__5981\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__6001\,
            I => \N__5978\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__5998\,
            I => \N__5975\
        );

    \I__1307\ : InMux
    port map (
            O => \N__5995\,
            I => \N__5972\
        );

    \I__1306\ : InMux
    port map (
            O => \N__5994\,
            I => \N__5964\
        );

    \I__1305\ : InMux
    port map (
            O => \N__5993\,
            I => \N__5964\
        );

    \I__1304\ : InMux
    port map (
            O => \N__5992\,
            I => \N__5964\
        );

    \I__1303\ : InMux
    port map (
            O => \N__5991\,
            I => \N__5961\
        );

    \I__1302\ : InMux
    port map (
            O => \N__5990\,
            I => \N__5954\
        );

    \I__1301\ : InMux
    port map (
            O => \N__5989\,
            I => \N__5954\
        );

    \I__1300\ : InMux
    port map (
            O => \N__5988\,
            I => \N__5954\
        );

    \I__1299\ : InMux
    port map (
            O => \N__5987\,
            I => \N__5951\
        );

    \I__1298\ : Span4Mux_v
    port map (
            O => \N__5984\,
            I => \N__5945\
        );

    \I__1297\ : Span4Mux_v
    port map (
            O => \N__5981\,
            I => \N__5945\
        );

    \I__1296\ : Span4Mux_v
    port map (
            O => \N__5978\,
            I => \N__5940\
        );

    \I__1295\ : Span4Mux_v
    port map (
            O => \N__5975\,
            I => \N__5940\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__5972\,
            I => \N__5937\
        );

    \I__1293\ : InMux
    port map (
            O => \N__5971\,
            I => \N__5934\
        );

    \I__1292\ : LocalMux
    port map (
            O => \N__5964\,
            I => \N__5924\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__5961\,
            I => \N__5924\
        );

    \I__1290\ : LocalMux
    port map (
            O => \N__5954\,
            I => \N__5924\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__5951\,
            I => \N__5924\
        );

    \I__1288\ : InMux
    port map (
            O => \N__5950\,
            I => \N__5921\
        );

    \I__1287\ : Sp12to4
    port map (
            O => \N__5945\,
            I => \N__5916\
        );

    \I__1286\ : Sp12to4
    port map (
            O => \N__5940\,
            I => \N__5916\
        );

    \I__1285\ : Span4Mux_h
    port map (
            O => \N__5937\,
            I => \N__5911\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__5934\,
            I => \N__5911\
        );

    \I__1283\ : InMux
    port map (
            O => \N__5933\,
            I => \N__5908\
        );

    \I__1282\ : Span4Mux_v
    port map (
            O => \N__5924\,
            I => \N__5903\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__5921\,
            I => \N__5903\
        );

    \I__1280\ : Odrv12
    port map (
            O => \N__5916\,
            I => columna_5
        );

    \I__1279\ : Odrv4
    port map (
            O => \N__5911\,
            I => columna_5
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__5908\,
            I => columna_5
        );

    \I__1277\ : Odrv4
    port map (
            O => \N__5903\,
            I => columna_5
        );

    \I__1276\ : InMux
    port map (
            O => \N__5894\,
            I => \N__5891\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__5891\,
            I => \N__5888\
        );

    \I__1274\ : Odrv12
    port map (
            O => \N__5888\,
            I => \generador.n1873\
        );

    \I__1273\ : CascadeMux
    port map (
            O => \N__5885\,
            I => \N__5882\
        );

    \I__1272\ : InMux
    port map (
            O => \N__5882\,
            I => \N__5879\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__5879\,
            I => \N__5872\
        );

    \I__1270\ : InMux
    port map (
            O => \N__5878\,
            I => \N__5866\
        );

    \I__1269\ : InMux
    port map (
            O => \N__5877\,
            I => \N__5866\
        );

    \I__1268\ : InMux
    port map (
            O => \N__5876\,
            I => \N__5861\
        );

    \I__1267\ : InMux
    port map (
            O => \N__5875\,
            I => \N__5861\
        );

    \I__1266\ : Span4Mux_h
    port map (
            O => \N__5872\,
            I => \N__5858\
        );

    \I__1265\ : InMux
    port map (
            O => \N__5871\,
            I => \N__5855\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__5866\,
            I => \N__5850\
        );

    \I__1263\ : LocalMux
    port map (
            O => \N__5861\,
            I => \N__5850\
        );

    \I__1262\ : Odrv4
    port map (
            O => \N__5858\,
            I => n14_adj_133
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__5855\,
            I => n14_adj_133
        );

    \I__1260\ : Odrv4
    port map (
            O => \N__5850\,
            I => n14_adj_133
        );

    \I__1259\ : CascadeMux
    port map (
            O => \N__5843\,
            I => \N__5840\
        );

    \I__1258\ : InMux
    port map (
            O => \N__5840\,
            I => \N__5835\
        );

    \I__1257\ : CascadeMux
    port map (
            O => \N__5839\,
            I => \N__5831\
        );

    \I__1256\ : InMux
    port map (
            O => \N__5838\,
            I => \N__5826\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__5835\,
            I => \N__5820\
        );

    \I__1254\ : InMux
    port map (
            O => \N__5834\,
            I => \N__5817\
        );

    \I__1253\ : InMux
    port map (
            O => \N__5831\,
            I => \N__5814\
        );

    \I__1252\ : InMux
    port map (
            O => \N__5830\,
            I => \N__5811\
        );

    \I__1251\ : CascadeMux
    port map (
            O => \N__5829\,
            I => \N__5807\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__5826\,
            I => \N__5804\
        );

    \I__1249\ : InMux
    port map (
            O => \N__5825\,
            I => \N__5801\
        );

    \I__1248\ : InMux
    port map (
            O => \N__5824\,
            I => \N__5796\
        );

    \I__1247\ : InMux
    port map (
            O => \N__5823\,
            I => \N__5796\
        );

    \I__1246\ : Span4Mux_h
    port map (
            O => \N__5820\,
            I => \N__5787\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__5817\,
            I => \N__5787\
        );

    \I__1244\ : LocalMux
    port map (
            O => \N__5814\,
            I => \N__5787\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__5811\,
            I => \N__5787\
        );

    \I__1242\ : InMux
    port map (
            O => \N__5810\,
            I => \N__5784\
        );

    \I__1241\ : InMux
    port map (
            O => \N__5807\,
            I => \N__5781\
        );

    \I__1240\ : Odrv4
    port map (
            O => \N__5804\,
            I => char_code_0
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__5801\,
            I => char_code_0
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__5796\,
            I => char_code_0
        );

    \I__1237\ : Odrv4
    port map (
            O => \N__5787\,
            I => char_code_0
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__5784\,
            I => char_code_0
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__5781\,
            I => char_code_0
        );

    \I__1234\ : CascadeMux
    port map (
            O => \N__5768\,
            I => \N__5765\
        );

    \I__1233\ : InMux
    port map (
            O => \N__5765\,
            I => \N__5754\
        );

    \I__1232\ : InMux
    port map (
            O => \N__5764\,
            I => \N__5754\
        );

    \I__1231\ : InMux
    port map (
            O => \N__5763\,
            I => \N__5750\
        );

    \I__1230\ : InMux
    port map (
            O => \N__5762\,
            I => \N__5745\
        );

    \I__1229\ : InMux
    port map (
            O => \N__5761\,
            I => \N__5745\
        );

    \I__1228\ : InMux
    port map (
            O => \N__5760\,
            I => \N__5742\
        );

    \I__1227\ : InMux
    port map (
            O => \N__5759\,
            I => \N__5739\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__5754\,
            I => \N__5736\
        );

    \I__1225\ : InMux
    port map (
            O => \N__5753\,
            I => \N__5733\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__5750\,
            I => n1166
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__5745\,
            I => n1166
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__5742\,
            I => n1166
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__5739\,
            I => n1166
        );

    \I__1220\ : Odrv4
    port map (
            O => \N__5736\,
            I => n1166
        );

    \I__1219\ : LocalMux
    port map (
            O => \N__5733\,
            I => n1166
        );

    \I__1218\ : InMux
    port map (
            O => \N__5720\,
            I => \N__5714\
        );

    \I__1217\ : InMux
    port map (
            O => \N__5719\,
            I => \N__5709\
        );

    \I__1216\ : InMux
    port map (
            O => \N__5718\,
            I => \N__5709\
        );

    \I__1215\ : InMux
    port map (
            O => \N__5717\,
            I => \N__5706\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__5714\,
            I => \N__5702\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__5709\,
            I => \N__5699\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__5706\,
            I => \N__5696\
        );

    \I__1211\ : CascadeMux
    port map (
            O => \N__5705\,
            I => \N__5689\
        );

    \I__1210\ : Span4Mux_v
    port map (
            O => \N__5702\,
            I => \N__5680\
        );

    \I__1209\ : Span4Mux_v
    port map (
            O => \N__5699\,
            I => \N__5680\
        );

    \I__1208\ : Span4Mux_v
    port map (
            O => \N__5696\,
            I => \N__5680\
        );

    \I__1207\ : InMux
    port map (
            O => \N__5695\,
            I => \N__5675\
        );

    \I__1206\ : InMux
    port map (
            O => \N__5694\,
            I => \N__5675\
        );

    \I__1205\ : InMux
    port map (
            O => \N__5693\,
            I => \N__5669\
        );

    \I__1204\ : InMux
    port map (
            O => \N__5692\,
            I => \N__5669\
        );

    \I__1203\ : InMux
    port map (
            O => \N__5689\,
            I => \N__5662\
        );

    \I__1202\ : InMux
    port map (
            O => \N__5688\,
            I => \N__5657\
        );

    \I__1201\ : InMux
    port map (
            O => \N__5687\,
            I => \N__5657\
        );

    \I__1200\ : Sp12to4
    port map (
            O => \N__5680\,
            I => \N__5652\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__5675\,
            I => \N__5652\
        );

    \I__1198\ : InMux
    port map (
            O => \N__5674\,
            I => \N__5649\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__5669\,
            I => \N__5646\
        );

    \I__1196\ : InMux
    port map (
            O => \N__5668\,
            I => \N__5641\
        );

    \I__1195\ : InMux
    port map (
            O => \N__5667\,
            I => \N__5641\
        );

    \I__1194\ : InMux
    port map (
            O => \N__5666\,
            I => \N__5638\
        );

    \I__1193\ : InMux
    port map (
            O => \N__5665\,
            I => \N__5635\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__5662\,
            I => n1212
        );

    \I__1191\ : LocalMux
    port map (
            O => \N__5657\,
            I => n1212
        );

    \I__1190\ : Odrv12
    port map (
            O => \N__5652\,
            I => n1212
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__5649\,
            I => n1212
        );

    \I__1188\ : Odrv4
    port map (
            O => \N__5646\,
            I => n1212
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__5641\,
            I => n1212
        );

    \I__1186\ : LocalMux
    port map (
            O => \N__5638\,
            I => n1212
        );

    \I__1185\ : LocalMux
    port map (
            O => \N__5635\,
            I => n1212
        );

    \I__1184\ : CascadeMux
    port map (
            O => \N__5618\,
            I => \tabla.n677_cascade_\
        );

    \I__1183\ : InMux
    port map (
            O => \N__5615\,
            I => \N__5612\
        );

    \I__1182\ : LocalMux
    port map (
            O => \N__5612\,
            I => \N__5609\
        );

    \I__1181\ : Odrv4
    port map (
            O => \N__5609\,
            I => \tabla.char_33\
        );

    \I__1180\ : InMux
    port map (
            O => \N__5606\,
            I => \N__5599\
        );

    \I__1179\ : InMux
    port map (
            O => \N__5605\,
            I => \N__5599\
        );

    \I__1178\ : InMux
    port map (
            O => \N__5604\,
            I => \N__5590\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__5599\,
            I => \N__5587\
        );

    \I__1176\ : InMux
    port map (
            O => \N__5598\,
            I => \N__5584\
        );

    \I__1175\ : InMux
    port map (
            O => \N__5597\,
            I => \N__5571\
        );

    \I__1174\ : InMux
    port map (
            O => \N__5596\,
            I => \N__5571\
        );

    \I__1173\ : InMux
    port map (
            O => \N__5595\,
            I => \N__5571\
        );

    \I__1172\ : InMux
    port map (
            O => \N__5594\,
            I => \N__5571\
        );

    \I__1171\ : InMux
    port map (
            O => \N__5593\,
            I => \N__5571\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__5590\,
            I => \N__5567\
        );

    \I__1169\ : Span4Mux_h
    port map (
            O => \N__5587\,
            I => \N__5562\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__5584\,
            I => \N__5562\
        );

    \I__1167\ : InMux
    port map (
            O => \N__5583\,
            I => \N__5559\
        );

    \I__1166\ : InMux
    port map (
            O => \N__5582\,
            I => \N__5554\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__5571\,
            I => \N__5551\
        );

    \I__1164\ : InMux
    port map (
            O => \N__5570\,
            I => \N__5548\
        );

    \I__1163\ : Span4Mux_v
    port map (
            O => \N__5567\,
            I => \N__5534\
        );

    \I__1162\ : Span4Mux_v
    port map (
            O => \N__5562\,
            I => \N__5529\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__5559\,
            I => \N__5529\
        );

    \I__1160\ : InMux
    port map (
            O => \N__5558\,
            I => \N__5524\
        );

    \I__1159\ : InMux
    port map (
            O => \N__5557\,
            I => \N__5524\
        );

    \I__1158\ : LocalMux
    port map (
            O => \N__5554\,
            I => \N__5517\
        );

    \I__1157\ : Span4Mux_h
    port map (
            O => \N__5551\,
            I => \N__5517\
        );

    \I__1156\ : LocalMux
    port map (
            O => \N__5548\,
            I => \N__5517\
        );

    \I__1155\ : InMux
    port map (
            O => \N__5547\,
            I => \N__5508\
        );

    \I__1154\ : InMux
    port map (
            O => \N__5546\,
            I => \N__5508\
        );

    \I__1153\ : InMux
    port map (
            O => \N__5545\,
            I => \N__5508\
        );

    \I__1152\ : InMux
    port map (
            O => \N__5544\,
            I => \N__5508\
        );

    \I__1151\ : InMux
    port map (
            O => \N__5543\,
            I => \N__5499\
        );

    \I__1150\ : InMux
    port map (
            O => \N__5542\,
            I => \N__5499\
        );

    \I__1149\ : InMux
    port map (
            O => \N__5541\,
            I => \N__5499\
        );

    \I__1148\ : InMux
    port map (
            O => \N__5540\,
            I => \N__5499\
        );

    \I__1147\ : InMux
    port map (
            O => \N__5539\,
            I => \N__5494\
        );

    \I__1146\ : InMux
    port map (
            O => \N__5538\,
            I => \N__5494\
        );

    \I__1145\ : InMux
    port map (
            O => \N__5537\,
            I => \N__5491\
        );

    \I__1144\ : Odrv4
    port map (
            O => \N__5534\,
            I => char_code_2
        );

    \I__1143\ : Odrv4
    port map (
            O => \N__5529\,
            I => char_code_2
        );

    \I__1142\ : LocalMux
    port map (
            O => \N__5524\,
            I => char_code_2
        );

    \I__1141\ : Odrv4
    port map (
            O => \N__5517\,
            I => char_code_2
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__5508\,
            I => char_code_2
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__5499\,
            I => char_code_2
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__5494\,
            I => char_code_2
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__5491\,
            I => char_code_2
        );

    \I__1136\ : CascadeMux
    port map (
            O => \N__5474\,
            I => \N__5463\
        );

    \I__1135\ : CascadeMux
    port map (
            O => \N__5473\,
            I => \N__5460\
        );

    \I__1134\ : CascadeMux
    port map (
            O => \N__5472\,
            I => \N__5457\
        );

    \I__1133\ : CascadeMux
    port map (
            O => \N__5471\,
            I => \N__5452\
        );

    \I__1132\ : CascadeMux
    port map (
            O => \N__5470\,
            I => \N__5449\
        );

    \I__1131\ : CascadeMux
    port map (
            O => \N__5469\,
            I => \N__5440\
        );

    \I__1130\ : CascadeMux
    port map (
            O => \N__5468\,
            I => \N__5435\
        );

    \I__1129\ : CascadeMux
    port map (
            O => \N__5467\,
            I => \N__5431\
        );

    \I__1128\ : InMux
    port map (
            O => \N__5466\,
            I => \N__5424\
        );

    \I__1127\ : InMux
    port map (
            O => \N__5463\,
            I => \N__5424\
        );

    \I__1126\ : InMux
    port map (
            O => \N__5460\,
            I => \N__5419\
        );

    \I__1125\ : InMux
    port map (
            O => \N__5457\,
            I => \N__5419\
        );

    \I__1124\ : InMux
    port map (
            O => \N__5456\,
            I => \N__5410\
        );

    \I__1123\ : InMux
    port map (
            O => \N__5455\,
            I => \N__5410\
        );

    \I__1122\ : InMux
    port map (
            O => \N__5452\,
            I => \N__5410\
        );

    \I__1121\ : InMux
    port map (
            O => \N__5449\,
            I => \N__5410\
        );

    \I__1120\ : InMux
    port map (
            O => \N__5448\,
            I => \N__5406\
        );

    \I__1119\ : InMux
    port map (
            O => \N__5447\,
            I => \N__5403\
        );

    \I__1118\ : InMux
    port map (
            O => \N__5446\,
            I => \N__5398\
        );

    \I__1117\ : InMux
    port map (
            O => \N__5445\,
            I => \N__5398\
        );

    \I__1116\ : InMux
    port map (
            O => \N__5444\,
            I => \N__5395\
        );

    \I__1115\ : InMux
    port map (
            O => \N__5443\,
            I => \N__5386\
        );

    \I__1114\ : InMux
    port map (
            O => \N__5440\,
            I => \N__5386\
        );

    \I__1113\ : InMux
    port map (
            O => \N__5439\,
            I => \N__5386\
        );

    \I__1112\ : InMux
    port map (
            O => \N__5438\,
            I => \N__5386\
        );

    \I__1111\ : InMux
    port map (
            O => \N__5435\,
            I => \N__5379\
        );

    \I__1110\ : InMux
    port map (
            O => \N__5434\,
            I => \N__5379\
        );

    \I__1109\ : InMux
    port map (
            O => \N__5431\,
            I => \N__5379\
        );

    \I__1108\ : InMux
    port map (
            O => \N__5430\,
            I => \N__5374\
        );

    \I__1107\ : InMux
    port map (
            O => \N__5429\,
            I => \N__5374\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__5424\,
            I => \N__5369\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__5419\,
            I => \N__5364\
        );

    \I__1104\ : LocalMux
    port map (
            O => \N__5410\,
            I => \N__5364\
        );

    \I__1103\ : InMux
    port map (
            O => \N__5409\,
            I => \N__5361\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__5406\,
            I => \N__5356\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__5403\,
            I => \N__5356\
        );

    \I__1100\ : LocalMux
    port map (
            O => \N__5398\,
            I => \N__5353\
        );

    \I__1099\ : LocalMux
    port map (
            O => \N__5395\,
            I => \N__5348\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__5386\,
            I => \N__5348\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__5379\,
            I => \N__5345\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__5374\,
            I => \N__5342\
        );

    \I__1095\ : InMux
    port map (
            O => \N__5373\,
            I => \N__5337\
        );

    \I__1094\ : InMux
    port map (
            O => \N__5372\,
            I => \N__5337\
        );

    \I__1093\ : Span4Mux_v
    port map (
            O => \N__5369\,
            I => \N__5332\
        );

    \I__1092\ : Span4Mux_v
    port map (
            O => \N__5364\,
            I => \N__5332\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__5361\,
            I => \N__5329\
        );

    \I__1090\ : Span4Mux_v
    port map (
            O => \N__5356\,
            I => \N__5316\
        );

    \I__1089\ : Span4Mux_h
    port map (
            O => \N__5353\,
            I => \N__5316\
        );

    \I__1088\ : Span4Mux_v
    port map (
            O => \N__5348\,
            I => \N__5316\
        );

    \I__1087\ : Span4Mux_v
    port map (
            O => \N__5345\,
            I => \N__5316\
        );

    \I__1086\ : Span4Mux_h
    port map (
            O => \N__5342\,
            I => \N__5316\
        );

    \I__1085\ : LocalMux
    port map (
            O => \N__5337\,
            I => \N__5316\
        );

    \I__1084\ : Odrv4
    port map (
            O => \N__5332\,
            I => char_code_1
        );

    \I__1083\ : Odrv4
    port map (
            O => \N__5329\,
            I => char_code_1
        );

    \I__1082\ : Odrv4
    port map (
            O => \N__5316\,
            I => char_code_1
        );

    \I__1081\ : InMux
    port map (
            O => \N__5309\,
            I => \N__5303\
        );

    \I__1080\ : InMux
    port map (
            O => \N__5308\,
            I => \N__5298\
        );

    \I__1079\ : InMux
    port map (
            O => \N__5307\,
            I => \N__5298\
        );

    \I__1078\ : InMux
    port map (
            O => \N__5306\,
            I => \N__5295\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__5303\,
            I => n891
        );

    \I__1076\ : LocalMux
    port map (
            O => \N__5298\,
            I => n891
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__5295\,
            I => n891
        );

    \I__1074\ : InMux
    port map (
            O => \N__5288\,
            I => \N__5277\
        );

    \I__1073\ : InMux
    port map (
            O => \N__5287\,
            I => \N__5277\
        );

    \I__1072\ : InMux
    port map (
            O => \N__5286\,
            I => \N__5274\
        );

    \I__1071\ : InMux
    port map (
            O => \N__5285\,
            I => \N__5269\
        );

    \I__1070\ : InMux
    port map (
            O => \N__5284\,
            I => \N__5269\
        );

    \I__1069\ : CascadeMux
    port map (
            O => \N__5283\,
            I => \N__5260\
        );

    \I__1068\ : CascadeMux
    port map (
            O => \N__5282\,
            I => \N__5242\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__5277\,
            I => \N__5239\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__5274\,
            I => \N__5234\
        );

    \I__1065\ : LocalMux
    port map (
            O => \N__5269\,
            I => \N__5234\
        );

    \I__1064\ : InMux
    port map (
            O => \N__5268\,
            I => \N__5227\
        );

    \I__1063\ : InMux
    port map (
            O => \N__5267\,
            I => \N__5227\
        );

    \I__1062\ : InMux
    port map (
            O => \N__5266\,
            I => \N__5227\
        );

    \I__1061\ : InMux
    port map (
            O => \N__5265\,
            I => \N__5221\
        );

    \I__1060\ : InMux
    port map (
            O => \N__5264\,
            I => \N__5221\
        );

    \I__1059\ : InMux
    port map (
            O => \N__5263\,
            I => \N__5214\
        );

    \I__1058\ : InMux
    port map (
            O => \N__5260\,
            I => \N__5214\
        );

    \I__1057\ : InMux
    port map (
            O => \N__5259\,
            I => \N__5214\
        );

    \I__1056\ : InMux
    port map (
            O => \N__5258\,
            I => \N__5209\
        );

    \I__1055\ : InMux
    port map (
            O => \N__5257\,
            I => \N__5209\
        );

    \I__1054\ : InMux
    port map (
            O => \N__5256\,
            I => \N__5206\
        );

    \I__1053\ : InMux
    port map (
            O => \N__5255\,
            I => \N__5203\
        );

    \I__1052\ : InMux
    port map (
            O => \N__5254\,
            I => \N__5196\
        );

    \I__1051\ : InMux
    port map (
            O => \N__5253\,
            I => \N__5196\
        );

    \I__1050\ : InMux
    port map (
            O => \N__5252\,
            I => \N__5196\
        );

    \I__1049\ : InMux
    port map (
            O => \N__5251\,
            I => \N__5187\
        );

    \I__1048\ : InMux
    port map (
            O => \N__5250\,
            I => \N__5187\
        );

    \I__1047\ : InMux
    port map (
            O => \N__5249\,
            I => \N__5187\
        );

    \I__1046\ : InMux
    port map (
            O => \N__5248\,
            I => \N__5187\
        );

    \I__1045\ : InMux
    port map (
            O => \N__5247\,
            I => \N__5182\
        );

    \I__1044\ : InMux
    port map (
            O => \N__5246\,
            I => \N__5182\
        );

    \I__1043\ : InMux
    port map (
            O => \N__5245\,
            I => \N__5177\
        );

    \I__1042\ : InMux
    port map (
            O => \N__5242\,
            I => \N__5177\
        );

    \I__1041\ : Span4Mux_v
    port map (
            O => \N__5239\,
            I => \N__5168\
        );

    \I__1040\ : Span4Mux_v
    port map (
            O => \N__5234\,
            I => \N__5168\
        );

    \I__1039\ : LocalMux
    port map (
            O => \N__5227\,
            I => \N__5168\
        );

    \I__1038\ : InMux
    port map (
            O => \N__5226\,
            I => \N__5165\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__5221\,
            I => \N__5158\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__5214\,
            I => \N__5158\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__5209\,
            I => \N__5158\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__5206\,
            I => \N__5149\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__5203\,
            I => \N__5149\
        );

    \I__1032\ : LocalMux
    port map (
            O => \N__5196\,
            I => \N__5149\
        );

    \I__1031\ : LocalMux
    port map (
            O => \N__5187\,
            I => \N__5149\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__5182\,
            I => \N__5144\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__5177\,
            I => \N__5144\
        );

    \I__1028\ : InMux
    port map (
            O => \N__5176\,
            I => \N__5141\
        );

    \I__1027\ : InMux
    port map (
            O => \N__5175\,
            I => \N__5138\
        );

    \I__1026\ : Span4Mux_h
    port map (
            O => \N__5168\,
            I => \N__5133\
        );

    \I__1025\ : LocalMux
    port map (
            O => \N__5165\,
            I => \N__5133\
        );

    \I__1024\ : Span4Mux_v
    port map (
            O => \N__5158\,
            I => \N__5122\
        );

    \I__1023\ : Span4Mux_v
    port map (
            O => \N__5149\,
            I => \N__5122\
        );

    \I__1022\ : Span4Mux_h
    port map (
            O => \N__5144\,
            I => \N__5122\
        );

    \I__1021\ : LocalMux
    port map (
            O => \N__5141\,
            I => \N__5122\
        );

    \I__1020\ : LocalMux
    port map (
            O => \N__5138\,
            I => \N__5122\
        );

    \I__1019\ : Odrv4
    port map (
            O => \N__5133\,
            I => char_code_3
        );

    \I__1018\ : Odrv4
    port map (
            O => \N__5122\,
            I => char_code_3
        );

    \I__1017\ : InMux
    port map (
            O => \N__5117\,
            I => \N__5114\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__5114\,
            I => \N__5110\
        );

    \I__1015\ : InMux
    port map (
            O => \N__5113\,
            I => \N__5107\
        );

    \I__1014\ : Odrv4
    port map (
            O => \N__5110\,
            I => \tabla.n876\
        );

    \I__1013\ : LocalMux
    port map (
            O => \N__5107\,
            I => \tabla.n876\
        );

    \I__1012\ : InMux
    port map (
            O => \N__5102\,
            I => \N__5099\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__5099\,
            I => \tabla.n1361\
        );

    \I__1010\ : InMux
    port map (
            O => \N__5096\,
            I => \N__5093\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__5093\,
            I => \tabla.char_38\
        );

    \I__1008\ : InMux
    port map (
            O => \N__5090\,
            I => \N__5087\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__5087\,
            I => \N__5083\
        );

    \I__1006\ : InMux
    port map (
            O => \N__5086\,
            I => \N__5080\
        );

    \I__1005\ : Odrv4
    port map (
            O => \N__5083\,
            I => char_36
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__5080\,
            I => char_36
        );

    \I__1003\ : InMux
    port map (
            O => \N__5075\,
            I => \N__5071\
        );

    \I__1002\ : InMux
    port map (
            O => \N__5074\,
            I => \N__5068\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__5071\,
            I => \N__5063\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__5068\,
            I => \N__5060\
        );

    \I__999\ : InMux
    port map (
            O => \N__5067\,
            I => \N__5055\
        );

    \I__998\ : InMux
    port map (
            O => \N__5066\,
            I => \N__5055\
        );

    \I__997\ : Odrv12
    port map (
            O => \N__5063\,
            I => char_17
        );

    \I__996\ : Odrv4
    port map (
            O => \N__5060\,
            I => char_17
        );

    \I__995\ : LocalMux
    port map (
            O => \N__5055\,
            I => char_17
        );

    \I__994\ : CascadeMux
    port map (
            O => \N__5048\,
            I => \N__5044\
        );

    \I__993\ : InMux
    port map (
            O => \N__5047\,
            I => \N__5020\
        );

    \I__992\ : InMux
    port map (
            O => \N__5044\,
            I => \N__5017\
        );

    \I__991\ : InMux
    port map (
            O => \N__5043\,
            I => \N__5012\
        );

    \I__990\ : InMux
    port map (
            O => \N__5042\,
            I => \N__5012\
        );

    \I__989\ : InMux
    port map (
            O => \N__5041\,
            I => \N__5005\
        );

    \I__988\ : InMux
    port map (
            O => \N__5040\,
            I => \N__5005\
        );

    \I__987\ : InMux
    port map (
            O => \N__5039\,
            I => \N__5005\
        );

    \I__986\ : InMux
    port map (
            O => \N__5038\,
            I => \N__5002\
        );

    \I__985\ : InMux
    port map (
            O => \N__5037\,
            I => \N__4997\
        );

    \I__984\ : InMux
    port map (
            O => \N__5036\,
            I => \N__4997\
        );

    \I__983\ : InMux
    port map (
            O => \N__5035\,
            I => \N__4988\
        );

    \I__982\ : InMux
    port map (
            O => \N__5034\,
            I => \N__4988\
        );

    \I__981\ : InMux
    port map (
            O => \N__5033\,
            I => \N__4988\
        );

    \I__980\ : InMux
    port map (
            O => \N__5032\,
            I => \N__4988\
        );

    \I__979\ : InMux
    port map (
            O => \N__5031\,
            I => \N__4985\
        );

    \I__978\ : InMux
    port map (
            O => \N__5030\,
            I => \N__4976\
        );

    \I__977\ : InMux
    port map (
            O => \N__5029\,
            I => \N__4976\
        );

    \I__976\ : InMux
    port map (
            O => \N__5028\,
            I => \N__4976\
        );

    \I__975\ : InMux
    port map (
            O => \N__5027\,
            I => \N__4973\
        );

    \I__974\ : InMux
    port map (
            O => \N__5026\,
            I => \N__4968\
        );

    \I__973\ : InMux
    port map (
            O => \N__5025\,
            I => \N__4968\
        );

    \I__972\ : InMux
    port map (
            O => \N__5024\,
            I => \N__4963\
        );

    \I__971\ : InMux
    port map (
            O => \N__5023\,
            I => \N__4963\
        );

    \I__970\ : LocalMux
    port map (
            O => \N__5020\,
            I => \N__4954\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__5017\,
            I => \N__4954\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__5012\,
            I => \N__4951\
        );

    \I__967\ : LocalMux
    port map (
            O => \N__5005\,
            I => \N__4948\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__5002\,
            I => \N__4939\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__4997\,
            I => \N__4939\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__4988\,
            I => \N__4939\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__4985\,
            I => \N__4939\
        );

    \I__962\ : InMux
    port map (
            O => \N__4984\,
            I => \N__4935\
        );

    \I__961\ : InMux
    port map (
            O => \N__4983\,
            I => \N__4932\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__4976\,
            I => \N__4923\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__4973\,
            I => \N__4923\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__4968\,
            I => \N__4923\
        );

    \I__957\ : LocalMux
    port map (
            O => \N__4963\,
            I => \N__4923\
        );

    \I__956\ : InMux
    port map (
            O => \N__4962\,
            I => \N__4916\
        );

    \I__955\ : InMux
    port map (
            O => \N__4961\,
            I => \N__4916\
        );

    \I__954\ : InMux
    port map (
            O => \N__4960\,
            I => \N__4916\
        );

    \I__953\ : InMux
    port map (
            O => \N__4959\,
            I => \N__4913\
        );

    \I__952\ : Span4Mux_v
    port map (
            O => \N__4954\,
            I => \N__4903\
        );

    \I__951\ : Span4Mux_v
    port map (
            O => \N__4951\,
            I => \N__4903\
        );

    \I__950\ : Span4Mux_v
    port map (
            O => \N__4948\,
            I => \N__4903\
        );

    \I__949\ : Span4Mux_v
    port map (
            O => \N__4939\,
            I => \N__4903\
        );

    \I__948\ : InMux
    port map (
            O => \N__4938\,
            I => \N__4900\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__4935\,
            I => \N__4894\
        );

    \I__946\ : LocalMux
    port map (
            O => \N__4932\,
            I => \N__4894\
        );

    \I__945\ : Span4Mux_v
    port map (
            O => \N__4923\,
            I => \N__4887\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__4916\,
            I => \N__4887\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__4913\,
            I => \N__4887\
        );

    \I__942\ : InMux
    port map (
            O => \N__4912\,
            I => \N__4884\
        );

    \I__941\ : Span4Mux_h
    port map (
            O => \N__4903\,
            I => \N__4881\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__4900\,
            I => \N__4878\
        );

    \I__939\ : InMux
    port map (
            O => \N__4899\,
            I => \N__4875\
        );

    \I__938\ : Span4Mux_v
    port map (
            O => \N__4894\,
            I => \N__4868\
        );

    \I__937\ : Span4Mux_h
    port map (
            O => \N__4887\,
            I => \N__4868\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__4884\,
            I => \N__4868\
        );

    \I__935\ : Odrv4
    port map (
            O => \N__4881\,
            I => columna_4
        );

    \I__934\ : Odrv4
    port map (
            O => \N__4878\,
            I => columna_4
        );

    \I__933\ : LocalMux
    port map (
            O => \N__4875\,
            I => columna_4
        );

    \I__932\ : Odrv4
    port map (
            O => \N__4868\,
            I => columna_4
        );

    \I__931\ : InMux
    port map (
            O => \N__4859\,
            I => \N__4856\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__4856\,
            I => \N__4853\
        );

    \I__929\ : Span4Mux_v
    port map (
            O => \N__4853\,
            I => \N__4850\
        );

    \I__928\ : Odrv4
    port map (
            O => \N__4850\,
            I => n24
        );

    \I__927\ : CascadeMux
    port map (
            O => \N__4847\,
            I => \n1347_cascade_\
        );

    \I__926\ : CascadeMux
    port map (
            O => \N__4844\,
            I => \N__4836\
        );

    \I__925\ : CascadeMux
    port map (
            O => \N__4843\,
            I => \N__4833\
        );

    \I__924\ : CascadeMux
    port map (
            O => \N__4842\,
            I => \N__4830\
        );

    \I__923\ : CascadeMux
    port map (
            O => \N__4841\,
            I => \N__4827\
        );

    \I__922\ : CascadeMux
    port map (
            O => \N__4840\,
            I => \N__4824\
        );

    \I__921\ : CascadeMux
    port map (
            O => \N__4839\,
            I => \N__4821\
        );

    \I__920\ : InMux
    port map (
            O => \N__4836\,
            I => \N__4815\
        );

    \I__919\ : InMux
    port map (
            O => \N__4833\,
            I => \N__4815\
        );

    \I__918\ : InMux
    port map (
            O => \N__4830\,
            I => \N__4810\
        );

    \I__917\ : InMux
    port map (
            O => \N__4827\,
            I => \N__4810\
        );

    \I__916\ : InMux
    port map (
            O => \N__4824\,
            I => \N__4798\
        );

    \I__915\ : InMux
    port map (
            O => \N__4821\,
            I => \N__4798\
        );

    \I__914\ : CascadeMux
    port map (
            O => \N__4820\,
            I => \N__4793\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__4815\,
            I => \N__4790\
        );

    \I__912\ : LocalMux
    port map (
            O => \N__4810\,
            I => \N__4787\
        );

    \I__911\ : InMux
    port map (
            O => \N__4809\,
            I => \N__4780\
        );

    \I__910\ : InMux
    port map (
            O => \N__4808\,
            I => \N__4780\
        );

    \I__909\ : InMux
    port map (
            O => \N__4807\,
            I => \N__4780\
        );

    \I__908\ : InMux
    port map (
            O => \N__4806\,
            I => \N__4777\
        );

    \I__907\ : InMux
    port map (
            O => \N__4805\,
            I => \N__4772\
        );

    \I__906\ : InMux
    port map (
            O => \N__4804\,
            I => \N__4772\
        );

    \I__905\ : InMux
    port map (
            O => \N__4803\,
            I => \N__4769\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__4798\,
            I => \N__4766\
        );

    \I__903\ : InMux
    port map (
            O => \N__4797\,
            I => \N__4761\
        );

    \I__902\ : InMux
    port map (
            O => \N__4796\,
            I => \N__4761\
        );

    \I__901\ : InMux
    port map (
            O => \N__4793\,
            I => \N__4758\
        );

    \I__900\ : Span4Mux_v
    port map (
            O => \N__4790\,
            I => \N__4752\
        );

    \I__899\ : Span4Mux_v
    port map (
            O => \N__4787\,
            I => \N__4752\
        );

    \I__898\ : LocalMux
    port map (
            O => \N__4780\,
            I => \N__4747\
        );

    \I__897\ : LocalMux
    port map (
            O => \N__4777\,
            I => \N__4747\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__4772\,
            I => \N__4742\
        );

    \I__895\ : LocalMux
    port map (
            O => \N__4769\,
            I => \N__4742\
        );

    \I__894\ : Span4Mux_v
    port map (
            O => \N__4766\,
            I => \N__4737\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__4761\,
            I => \N__4737\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__4758\,
            I => \N__4734\
        );

    \I__891\ : InMux
    port map (
            O => \N__4757\,
            I => \N__4731\
        );

    \I__890\ : Span4Mux_h
    port map (
            O => \N__4752\,
            I => \N__4726\
        );

    \I__889\ : Span4Mux_v
    port map (
            O => \N__4747\,
            I => \N__4726\
        );

    \I__888\ : Odrv12
    port map (
            O => \N__4742\,
            I => columna_8
        );

    \I__887\ : Odrv4
    port map (
            O => \N__4737\,
            I => columna_8
        );

    \I__886\ : Odrv4
    port map (
            O => \N__4734\,
            I => columna_8
        );

    \I__885\ : LocalMux
    port map (
            O => \N__4731\,
            I => columna_8
        );

    \I__884\ : Odrv4
    port map (
            O => \N__4726\,
            I => columna_8
        );

    \I__883\ : InMux
    port map (
            O => \N__4715\,
            I => \N__4702\
        );

    \I__882\ : InMux
    port map (
            O => \N__4714\,
            I => \N__4702\
        );

    \I__881\ : InMux
    port map (
            O => \N__4713\,
            I => \N__4691\
        );

    \I__880\ : InMux
    port map (
            O => \N__4712\,
            I => \N__4691\
        );

    \I__879\ : InMux
    port map (
            O => \N__4711\,
            I => \N__4686\
        );

    \I__878\ : InMux
    port map (
            O => \N__4710\,
            I => \N__4686\
        );

    \I__877\ : InMux
    port map (
            O => \N__4709\,
            I => \N__4679\
        );

    \I__876\ : InMux
    port map (
            O => \N__4708\,
            I => \N__4679\
        );

    \I__875\ : InMux
    port map (
            O => \N__4707\,
            I => \N__4679\
        );

    \I__874\ : LocalMux
    port map (
            O => \N__4702\,
            I => \N__4674\
        );

    \I__873\ : InMux
    port map (
            O => \N__4701\,
            I => \N__4669\
        );

    \I__872\ : InMux
    port map (
            O => \N__4700\,
            I => \N__4669\
        );

    \I__871\ : InMux
    port map (
            O => \N__4699\,
            I => \N__4662\
        );

    \I__870\ : InMux
    port map (
            O => \N__4698\,
            I => \N__4662\
        );

    \I__869\ : InMux
    port map (
            O => \N__4697\,
            I => \N__4662\
        );

    \I__868\ : InMux
    port map (
            O => \N__4696\,
            I => \N__4659\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__4691\,
            I => \N__4656\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__4686\,
            I => \N__4653\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__4679\,
            I => \N__4650\
        );

    \I__864\ : InMux
    port map (
            O => \N__4678\,
            I => \N__4647\
        );

    \I__863\ : InMux
    port map (
            O => \N__4677\,
            I => \N__4644\
        );

    \I__862\ : Span4Mux_v
    port map (
            O => \N__4674\,
            I => \N__4638\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__4669\,
            I => \N__4638\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__4662\,
            I => \N__4633\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__4659\,
            I => \N__4633\
        );

    \I__858\ : Span12Mux_h
    port map (
            O => \N__4656\,
            I => \N__4630\
        );

    \I__857\ : Span4Mux_v
    port map (
            O => \N__4653\,
            I => \N__4623\
        );

    \I__856\ : Span4Mux_v
    port map (
            O => \N__4650\,
            I => \N__4623\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__4647\,
            I => \N__4623\
        );

    \I__854\ : LocalMux
    port map (
            O => \N__4644\,
            I => \N__4620\
        );

    \I__853\ : InMux
    port map (
            O => \N__4643\,
            I => \N__4617\
        );

    \I__852\ : Span4Mux_h
    port map (
            O => \N__4638\,
            I => \N__4612\
        );

    \I__851\ : Span4Mux_v
    port map (
            O => \N__4633\,
            I => \N__4612\
        );

    \I__850\ : Odrv12
    port map (
            O => \N__4630\,
            I => columna_9
        );

    \I__849\ : Odrv4
    port map (
            O => \N__4623\,
            I => columna_9
        );

    \I__848\ : Odrv4
    port map (
            O => \N__4620\,
            I => columna_9
        );

    \I__847\ : LocalMux
    port map (
            O => \N__4617\,
            I => columna_9
        );

    \I__846\ : Odrv4
    port map (
            O => \N__4612\,
            I => columna_9
        );

    \I__845\ : InMux
    port map (
            O => \N__4601\,
            I => \N__4598\
        );

    \I__844\ : LocalMux
    port map (
            O => \N__4598\,
            I => \tabla.n1930\
        );

    \I__843\ : CascadeMux
    port map (
            O => \N__4595\,
            I => \N__4592\
        );

    \I__842\ : InMux
    port map (
            O => \N__4592\,
            I => \N__4587\
        );

    \I__841\ : InMux
    port map (
            O => \N__4591\,
            I => \N__4584\
        );

    \I__840\ : InMux
    port map (
            O => \N__4590\,
            I => \N__4579\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__4587\,
            I => \N__4576\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__4584\,
            I => \N__4573\
        );

    \I__837\ : InMux
    port map (
            O => \N__4583\,
            I => \N__4568\
        );

    \I__836\ : InMux
    port map (
            O => \N__4582\,
            I => \N__4568\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__4579\,
            I => \tabla.n1349\
        );

    \I__834\ : Odrv4
    port map (
            O => \N__4576\,
            I => \tabla.n1349\
        );

    \I__833\ : Odrv12
    port map (
            O => \N__4573\,
            I => \tabla.n1349\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__4568\,
            I => \tabla.n1349\
        );

    \I__831\ : CascadeMux
    port map (
            O => \N__4559\,
            I => \tabla.n1930_cascade_\
        );

    \I__830\ : InMux
    port map (
            O => \N__4556\,
            I => \N__4553\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__4553\,
            I => n1994
        );

    \I__828\ : InMux
    port map (
            O => \N__4550\,
            I => \N__4547\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__4547\,
            I => \tabla.n7_adj_127\
        );

    \I__826\ : InMux
    port map (
            O => \N__4544\,
            I => \N__4540\
        );

    \I__825\ : InMux
    port map (
            O => \N__4543\,
            I => \N__4537\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__4540\,
            I => char_19
        );

    \I__823\ : LocalMux
    port map (
            O => \N__4537\,
            I => char_19
        );

    \I__822\ : CascadeMux
    port map (
            O => \N__4532\,
            I => \N__4526\
        );

    \I__821\ : InMux
    port map (
            O => \N__4531\,
            I => \N__4517\
        );

    \I__820\ : InMux
    port map (
            O => \N__4530\,
            I => \N__4514\
        );

    \I__819\ : InMux
    port map (
            O => \N__4529\,
            I => \N__4511\
        );

    \I__818\ : InMux
    port map (
            O => \N__4526\,
            I => \N__4502\
        );

    \I__817\ : InMux
    port map (
            O => \N__4525\,
            I => \N__4502\
        );

    \I__816\ : InMux
    port map (
            O => \N__4524\,
            I => \N__4502\
        );

    \I__815\ : InMux
    port map (
            O => \N__4523\,
            I => \N__4502\
        );

    \I__814\ : InMux
    port map (
            O => \N__4522\,
            I => \N__4499\
        );

    \I__813\ : InMux
    port map (
            O => \N__4521\,
            I => \N__4494\
        );

    \I__812\ : InMux
    port map (
            O => \N__4520\,
            I => \N__4494\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__4517\,
            I => \N__4485\
        );

    \I__810\ : LocalMux
    port map (
            O => \N__4514\,
            I => \N__4485\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__4511\,
            I => \N__4485\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__4502\,
            I => \N__4482\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__4499\,
            I => \N__4477\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__4494\,
            I => \N__4477\
        );

    \I__805\ : InMux
    port map (
            O => \N__4493\,
            I => \N__4473\
        );

    \I__804\ : InMux
    port map (
            O => \N__4492\,
            I => \N__4470\
        );

    \I__803\ : Span4Mux_v
    port map (
            O => \N__4485\,
            I => \N__4465\
        );

    \I__802\ : Span4Mux_v
    port map (
            O => \N__4482\,
            I => \N__4460\
        );

    \I__801\ : Span4Mux_h
    port map (
            O => \N__4477\,
            I => \N__4460\
        );

    \I__800\ : InMux
    port map (
            O => \N__4476\,
            I => \N__4457\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__4473\,
            I => \N__4452\
        );

    \I__798\ : LocalMux
    port map (
            O => \N__4470\,
            I => \N__4452\
        );

    \I__797\ : InMux
    port map (
            O => \N__4469\,
            I => \N__4449\
        );

    \I__796\ : InMux
    port map (
            O => \N__4468\,
            I => \N__4446\
        );

    \I__795\ : Span4Mux_h
    port map (
            O => \N__4465\,
            I => \N__4443\
        );

    \I__794\ : Span4Mux_h
    port map (
            O => \N__4460\,
            I => \N__4438\
        );

    \I__793\ : LocalMux
    port map (
            O => \N__4457\,
            I => \N__4438\
        );

    \I__792\ : Span4Mux_v
    port map (
            O => \N__4452\,
            I => \N__4431\
        );

    \I__791\ : LocalMux
    port map (
            O => \N__4449\,
            I => \N__4431\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__4446\,
            I => \N__4431\
        );

    \I__789\ : Odrv4
    port map (
            O => \N__4443\,
            I => columna_6
        );

    \I__788\ : Odrv4
    port map (
            O => \N__4438\,
            I => columna_6
        );

    \I__787\ : Odrv4
    port map (
            O => \N__4431\,
            I => columna_6
        );

    \I__786\ : InMux
    port map (
            O => \N__4424\,
            I => \N__4421\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__4421\,
            I => \N__4418\
        );

    \I__784\ : Odrv12
    port map (
            O => \N__4418\,
            I => \generador.n1976\
        );

    \I__783\ : CascadeMux
    port map (
            O => \N__4415\,
            I => \n17_cascade_\
        );

    \I__782\ : InMux
    port map (
            O => \N__4412\,
            I => \N__4409\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__4409\,
            I => \N__4406\
        );

    \I__780\ : Span4Mux_v
    port map (
            O => \N__4406\,
            I => \N__4403\
        );

    \I__779\ : Odrv4
    port map (
            O => \N__4403\,
            I => \generador.n1979\
        );

    \I__778\ : InMux
    port map (
            O => \N__4400\,
            I => \N__4396\
        );

    \I__777\ : InMux
    port map (
            O => \N__4399\,
            I => \N__4393\
        );

    \I__776\ : LocalMux
    port map (
            O => \N__4396\,
            I => \N__4385\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__4393\,
            I => \N__4385\
        );

    \I__774\ : InMux
    port map (
            O => \N__4392\,
            I => \N__4382\
        );

    \I__773\ : InMux
    port map (
            O => \N__4391\,
            I => \N__4377\
        );

    \I__772\ : InMux
    port map (
            O => \N__4390\,
            I => \N__4377\
        );

    \I__771\ : Odrv4
    port map (
            O => \N__4385\,
            I => \tabla.n1397\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__4382\,
            I => \tabla.n1397\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__4377\,
            I => \tabla.n1397\
        );

    \I__768\ : InMux
    port map (
            O => \N__4370\,
            I => \N__4367\
        );

    \I__767\ : LocalMux
    port map (
            O => \N__4367\,
            I => n16
        );

    \I__766\ : CascadeMux
    port map (
            O => \N__4364\,
            I => \N__4360\
        );

    \I__765\ : InMux
    port map (
            O => \N__4363\,
            I => \N__4355\
        );

    \I__764\ : InMux
    port map (
            O => \N__4360\,
            I => \N__4355\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__4355\,
            I => \N__4351\
        );

    \I__762\ : InMux
    port map (
            O => \N__4354\,
            I => \N__4348\
        );

    \I__761\ : Odrv4
    port map (
            O => \N__4351\,
            I => n1220
        );

    \I__760\ : LocalMux
    port map (
            O => \N__4348\,
            I => n1220
        );

    \I__759\ : CascadeMux
    port map (
            O => \N__4343\,
            I => \char_22_cascade_\
        );

    \I__758\ : CascadeMux
    port map (
            O => \N__4340\,
            I => \n19_cascade_\
        );

    \I__757\ : CascadeMux
    port map (
            O => \N__4337\,
            I => \tabla.n14_cascade_\
        );

    \I__756\ : InMux
    port map (
            O => \N__4334\,
            I => \N__4331\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__4331\,
            I => char_20
        );

    \I__754\ : InMux
    port map (
            O => \N__4328\,
            I => \N__4325\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__4325\,
            I => char_22
        );

    \I__752\ : InMux
    port map (
            O => \N__4322\,
            I => \N__4319\
        );

    \I__751\ : LocalMux
    port map (
            O => \N__4319\,
            I => n20
        );

    \I__750\ : InMux
    port map (
            O => \N__4316\,
            I => \N__4308\
        );

    \I__749\ : InMux
    port map (
            O => \N__4315\,
            I => \N__4308\
        );

    \I__748\ : InMux
    port map (
            O => \N__4314\,
            I => \N__4303\
        );

    \I__747\ : InMux
    port map (
            O => \N__4313\,
            I => \N__4303\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__4308\,
            I => n1385
        );

    \I__745\ : LocalMux
    port map (
            O => \N__4303\,
            I => n1385
        );

    \I__744\ : InMux
    port map (
            O => \N__4298\,
            I => \N__4294\
        );

    \I__743\ : InMux
    port map (
            O => \N__4297\,
            I => \N__4291\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__4294\,
            I => n1405
        );

    \I__741\ : LocalMux
    port map (
            O => \N__4291\,
            I => n1405
        );

    \I__740\ : InMux
    port map (
            O => \N__4286\,
            I => \N__4283\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__4283\,
            I => \tabla.n7\
        );

    \I__738\ : InMux
    port map (
            O => \N__4280\,
            I => \N__4276\
        );

    \I__737\ : CascadeMux
    port map (
            O => \N__4279\,
            I => \N__4272\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__4276\,
            I => \N__4267\
        );

    \I__735\ : InMux
    port map (
            O => \N__4275\,
            I => \N__4264\
        );

    \I__734\ : InMux
    port map (
            O => \N__4272\,
            I => \N__4261\
        );

    \I__733\ : InMux
    port map (
            O => \N__4271\,
            I => \N__4256\
        );

    \I__732\ : InMux
    port map (
            O => \N__4270\,
            I => \N__4256\
        );

    \I__731\ : Odrv4
    port map (
            O => \N__4267\,
            I => n1347
        );

    \I__730\ : LocalMux
    port map (
            O => \N__4264\,
            I => n1347
        );

    \I__729\ : LocalMux
    port map (
            O => \N__4261\,
            I => n1347
        );

    \I__728\ : LocalMux
    port map (
            O => \N__4256\,
            I => n1347
        );

    \I__727\ : CascadeMux
    port map (
            O => \N__4247\,
            I => \generador.n1608_cascade_\
        );

    \I__726\ : InMux
    port map (
            O => \N__4244\,
            I => \N__4241\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__4241\,
            I => \generador.n1008\
        );

    \I__724\ : CascadeMux
    port map (
            O => \N__4238\,
            I => \n1934_cascade_\
        );

    \I__723\ : InMux
    port map (
            O => \N__4235\,
            I => \N__4232\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__4232\,
            I => \N__4229\
        );

    \I__721\ : Odrv4
    port map (
            O => \N__4229\,
            I => \generador.n1021\
        );

    \I__720\ : InMux
    port map (
            O => \N__4226\,
            I => \N__4223\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__4223\,
            I => n51
        );

    \I__718\ : InMux
    port map (
            O => \N__4220\,
            I => \N__4217\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__4217\,
            I => \N__4214\
        );

    \I__716\ : Span4Mux_v
    port map (
            O => \N__4214\,
            I => \N__4209\
        );

    \I__715\ : InMux
    port map (
            O => \N__4213\,
            I => \N__4206\
        );

    \I__714\ : InMux
    port map (
            O => \N__4212\,
            I => \N__4203\
        );

    \I__713\ : Odrv4
    port map (
            O => \N__4209\,
            I => char_61
        );

    \I__712\ : LocalMux
    port map (
            O => \N__4206\,
            I => char_61
        );

    \I__711\ : LocalMux
    port map (
            O => \N__4203\,
            I => char_61
        );

    \I__710\ : CascadeMux
    port map (
            O => \N__4196\,
            I => \tabla.n1361_cascade_\
        );

    \I__709\ : CascadeMux
    port map (
            O => \N__4193\,
            I => \n1415_cascade_\
        );

    \I__708\ : InMux
    port map (
            O => \N__4190\,
            I => \N__4187\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__4187\,
            I => n1420
        );

    \I__706\ : CascadeMux
    port map (
            O => \N__4184\,
            I => \n1166_cascade_\
        );

    \I__705\ : CascadeMux
    port map (
            O => \N__4181\,
            I => \tabla.n7_adj_122_cascade_\
        );

    \I__704\ : InMux
    port map (
            O => \N__4178\,
            I => \N__4175\
        );

    \I__703\ : LocalMux
    port map (
            O => \N__4175\,
            I => \generador.n1019\
        );

    \I__702\ : InMux
    port map (
            O => \N__4172\,
            I => \N__4169\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__4169\,
            I => n5
        );

    \I__700\ : CascadeMux
    port map (
            O => \N__4166\,
            I => \N__4163\
        );

    \I__699\ : InMux
    port map (
            O => \N__4163\,
            I => \N__4160\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__4160\,
            I => n4
        );

    \I__697\ : CascadeMux
    port map (
            O => \N__4157\,
            I => \N__4152\
        );

    \I__696\ : CascadeMux
    port map (
            O => \N__4156\,
            I => \N__4144\
        );

    \I__695\ : InMux
    port map (
            O => \N__4155\,
            I => \N__4139\
        );

    \I__694\ : InMux
    port map (
            O => \N__4152\,
            I => \N__4139\
        );

    \I__693\ : InMux
    port map (
            O => \N__4151\,
            I => \N__4132\
        );

    \I__692\ : InMux
    port map (
            O => \N__4150\,
            I => \N__4132\
        );

    \I__691\ : InMux
    port map (
            O => \N__4149\,
            I => \N__4132\
        );

    \I__690\ : InMux
    port map (
            O => \N__4148\,
            I => \N__4129\
        );

    \I__689\ : InMux
    port map (
            O => \N__4147\,
            I => \N__4126\
        );

    \I__688\ : InMux
    port map (
            O => \N__4144\,
            I => \N__4123\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__4139\,
            I => n7_adj_137
        );

    \I__686\ : LocalMux
    port map (
            O => \N__4132\,
            I => n7_adj_137
        );

    \I__685\ : LocalMux
    port map (
            O => \N__4129\,
            I => n7_adj_137
        );

    \I__684\ : LocalMux
    port map (
            O => \N__4126\,
            I => n7_adj_137
        );

    \I__683\ : LocalMux
    port map (
            O => \N__4123\,
            I => n7_adj_137
        );

    \I__682\ : InMux
    port map (
            O => \N__4112\,
            I => \N__4106\
        );

    \I__681\ : InMux
    port map (
            O => \N__4111\,
            I => \N__4106\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__4106\,
            I => \N__4102\
        );

    \I__679\ : InMux
    port map (
            O => \N__4105\,
            I => \N__4099\
        );

    \I__678\ : Odrv4
    port map (
            O => \N__4102\,
            I => char_60
        );

    \I__677\ : LocalMux
    port map (
            O => \N__4099\,
            I => char_60
        );

    \I__676\ : InMux
    port map (
            O => \N__4094\,
            I => \N__4091\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__4091\,
            I => \N__4088\
        );

    \I__674\ : Odrv4
    port map (
            O => \N__4088\,
            I => n2
        );

    \I__673\ : InMux
    port map (
            O => \N__4085\,
            I => \N__4082\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__4082\,
            I => \generador.n1982\
        );

    \I__671\ : InMux
    port map (
            O => \N__4079\,
            I => \N__4076\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__4076\,
            I => \N__4073\
        );

    \I__669\ : Odrv12
    port map (
            O => \N__4073\,
            I => \generador.n1985\
        );

    \I__668\ : InMux
    port map (
            O => \N__4070\,
            I => \N__4067\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__4067\,
            I => \tabla.char_1\
        );

    \I__666\ : CascadeMux
    port map (
            O => \N__4064\,
            I => \N__4061\
        );

    \I__665\ : InMux
    port map (
            O => \N__4061\,
            I => \N__4058\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__4058\,
            I => n1
        );

    \I__663\ : CascadeMux
    port map (
            O => \N__4055\,
            I => \n7_cascade_\
        );

    \I__662\ : CascadeMux
    port map (
            O => \N__4052\,
            I => \n1012_cascade_\
        );

    \I__661\ : InMux
    port map (
            O => \N__4049\,
            I => \N__4046\
        );

    \I__660\ : LocalMux
    port map (
            O => \N__4046\,
            I => \generador.n1013\
        );

    \I__659\ : InMux
    port map (
            O => \N__4043\,
            I => \N__4040\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__4040\,
            I => n7
        );

    \I__657\ : CascadeMux
    port map (
            O => \N__4037\,
            I => \char_5_cascade_\
        );

    \I__656\ : InMux
    port map (
            O => \N__4034\,
            I => \N__4029\
        );

    \I__655\ : InMux
    port map (
            O => \N__4033\,
            I => \N__4024\
        );

    \I__654\ : InMux
    port map (
            O => \N__4032\,
            I => \N__4024\
        );

    \I__653\ : LocalMux
    port map (
            O => \N__4029\,
            I => char_11
        );

    \I__652\ : LocalMux
    port map (
            O => \N__4024\,
            I => char_11
        );

    \I__651\ : CascadeMux
    port map (
            O => \N__4019\,
            I => \char_code_0_cascade_\
        );

    \I__650\ : InMux
    port map (
            O => \N__4016\,
            I => \N__4013\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__4013\,
            I => \N__4010\
        );

    \I__648\ : Odrv4
    port map (
            O => \N__4010\,
            I => n1382
        );

    \I__647\ : CascadeMux
    port map (
            O => \N__4007\,
            I => \generador.n2006_cascade_\
        );

    \I__646\ : InMux
    port map (
            O => \N__4004\,
            I => \N__4001\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__4001\,
            I => \generador.n1847\
        );

    \I__644\ : CascadeMux
    port map (
            O => \N__3998\,
            I => \char_13_cascade_\
        );

    \I__643\ : CascadeMux
    port map (
            O => \N__3995\,
            I => \n11_cascade_\
        );

    \I__642\ : InMux
    port map (
            O => \N__3992\,
            I => \N__3989\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__3989\,
            I => \generador.n1988\
        );

    \I__640\ : CascadeMux
    port map (
            O => \N__3986\,
            I => \n1410_cascade_\
        );

    \I__639\ : InMux
    port map (
            O => \N__3983\,
            I => \N__3980\
        );

    \I__638\ : LocalMux
    port map (
            O => \N__3980\,
            I => \N__3977\
        );

    \I__637\ : Span4Mux_h
    port map (
            O => \N__3977\,
            I => \N__3974\
        );

    \I__636\ : Odrv4
    port map (
            O => \N__3974\,
            I => \generador.n1991\
        );

    \I__635\ : CascadeMux
    port map (
            O => \N__3971\,
            I => \tabla.char_14_cascade_\
        );

    \I__634\ : InMux
    port map (
            O => \N__3968\,
            I => \N__3965\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__3965\,
            I => n12
        );

    \I__632\ : InMux
    port map (
            O => \N__3962\,
            I => \N__3959\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__3959\,
            I => \generador.n1852\
        );

    \I__630\ : InMux
    port map (
            O => \N__3956\,
            I => \N__3953\
        );

    \I__629\ : LocalMux
    port map (
            O => \N__3953\,
            I => char_43
        );

    \I__628\ : CascadeMux
    port map (
            O => \N__3950\,
            I => \tabla.n728_cascade_\
        );

    \I__627\ : CascadeMux
    port map (
            O => \N__3947\,
            I => \N__3944\
        );

    \I__626\ : InMux
    port map (
            O => \N__3944\,
            I => \N__3941\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__3941\,
            I => char_50
        );

    \I__624\ : InMux
    port map (
            O => \N__3938\,
            I => \N__3935\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__3935\,
            I => n1952
        );

    \I__622\ : InMux
    port map (
            O => \N__3932\,
            I => \N__3929\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__3929\,
            I => n58
        );

    \I__620\ : CascadeMux
    port map (
            O => \N__3926\,
            I => \n57_cascade_\
        );

    \I__619\ : InMux
    port map (
            O => \N__3923\,
            I => \N__3920\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__3920\,
            I => \N__3917\
        );

    \I__617\ : Odrv4
    port map (
            O => \N__3917\,
            I => n54
        );

    \I__616\ : InMux
    port map (
            O => \N__3914\,
            I => \N__3911\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__3911\,
            I => n55
        );

    \I__614\ : CascadeMux
    port map (
            O => \N__3908\,
            I => \generador.n1964_cascade_\
        );

    \I__613\ : InMux
    port map (
            O => \N__3905\,
            I => \N__3902\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__3902\,
            I => \generador.n1967\
        );

    \I__611\ : InMux
    port map (
            O => \N__3899\,
            I => \N__3895\
        );

    \I__610\ : InMux
    port map (
            O => \N__3898\,
            I => \N__3892\
        );

    \I__609\ : LocalMux
    port map (
            O => \N__3895\,
            I => n1389
        );

    \I__608\ : LocalMux
    port map (
            O => \N__3892\,
            I => n1389
        );

    \I__607\ : InMux
    port map (
            O => \N__3887\,
            I => \N__3884\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__3884\,
            I => n42
        );

    \I__605\ : InMux
    port map (
            O => \N__3881\,
            I => \N__3877\
        );

    \I__604\ : InMux
    port map (
            O => \N__3880\,
            I => \N__3874\
        );

    \I__603\ : LocalMux
    port map (
            O => \N__3877\,
            I => \sincronismo.n1210\
        );

    \I__602\ : LocalMux
    port map (
            O => \N__3874\,
            I => \sincronismo.n1210\
        );

    \I__601\ : InMux
    port map (
            O => \N__3869\,
            I => \N__3865\
        );

    \I__600\ : InMux
    port map (
            O => \N__3868\,
            I => \N__3862\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__3865\,
            I => \sincronismo.n1932\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__3862\,
            I => \sincronismo.n1932\
        );

    \I__597\ : CascadeMux
    port map (
            O => \N__3857\,
            I => \n1212_cascade_\
        );

    \I__596\ : InMux
    port map (
            O => \N__3854\,
            I => \N__3851\
        );

    \I__595\ : LocalMux
    port map (
            O => \N__3851\,
            I => \tabla.n7_adj_124\
        );

    \I__594\ : InMux
    port map (
            O => \N__3848\,
            I => \N__3845\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__3845\,
            I => \sincronismo.n15_adj_117\
        );

    \I__592\ : CascadeMux
    port map (
            O => \N__3842\,
            I => \N__3839\
        );

    \I__591\ : InMux
    port map (
            O => \N__3839\,
            I => \N__3836\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__3836\,
            I => \sincronismo.n16\
        );

    \I__589\ : CascadeMux
    port map (
            O => \N__3833\,
            I => \N__3828\
        );

    \I__588\ : CascadeMux
    port map (
            O => \N__3832\,
            I => \N__3824\
        );

    \I__587\ : InMux
    port map (
            O => \N__3831\,
            I => \N__3819\
        );

    \I__586\ : InMux
    port map (
            O => \N__3828\,
            I => \N__3816\
        );

    \I__585\ : InMux
    port map (
            O => \N__3827\,
            I => \N__3812\
        );

    \I__584\ : InMux
    port map (
            O => \N__3824\,
            I => \N__3805\
        );

    \I__583\ : InMux
    port map (
            O => \N__3823\,
            I => \N__3805\
        );

    \I__582\ : InMux
    port map (
            O => \N__3822\,
            I => \N__3805\
        );

    \I__581\ : LocalMux
    port map (
            O => \N__3819\,
            I => \N__3798\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__3816\,
            I => \N__3798\
        );

    \I__579\ : InMux
    port map (
            O => \N__3815\,
            I => \N__3795\
        );

    \I__578\ : LocalMux
    port map (
            O => \N__3812\,
            I => \N__3792\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__3805\,
            I => \N__3789\
        );

    \I__576\ : InMux
    port map (
            O => \N__3804\,
            I => \N__3786\
        );

    \I__575\ : InMux
    port map (
            O => \N__3803\,
            I => \N__3783\
        );

    \I__574\ : Span4Mux_h
    port map (
            O => \N__3798\,
            I => \N__3780\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__3795\,
            I => \N__3777\
        );

    \I__572\ : Span4Mux_v
    port map (
            O => \N__3792\,
            I => \N__3768\
        );

    \I__571\ : Span4Mux_v
    port map (
            O => \N__3789\,
            I => \N__3768\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__3786\,
            I => \N__3768\
        );

    \I__569\ : LocalMux
    port map (
            O => \N__3783\,
            I => \N__3768\
        );

    \I__568\ : Odrv4
    port map (
            O => \N__3780\,
            I => columna_7
        );

    \I__567\ : Odrv4
    port map (
            O => \N__3777\,
            I => columna_7
        );

    \I__566\ : Odrv4
    port map (
            O => \N__3768\,
            I => columna_7
        );

    \I__565\ : InMux
    port map (
            O => \N__3761\,
            I => \N__3758\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__3758\,
            I => \tabla.n7_adj_129\
        );

    \I__563\ : CascadeMux
    port map (
            O => \N__3755\,
            I => \tabla.n7_adj_129_cascade_\
        );

    \I__562\ : InMux
    port map (
            O => \N__3752\,
            I => \N__3749\
        );

    \I__561\ : LocalMux
    port map (
            O => \N__3749\,
            I => \tabla.char_49\
        );

    \I__560\ : CascadeMux
    port map (
            O => \N__3746\,
            I => \tabla.n7_adj_128_cascade_\
        );

    \I__559\ : CascadeMux
    port map (
            O => \N__3743\,
            I => \N__3739\
        );

    \I__558\ : InMux
    port map (
            O => \N__3742\,
            I => \N__3734\
        );

    \I__557\ : InMux
    port map (
            O => \N__3739\,
            I => \N__3734\
        );

    \I__556\ : LocalMux
    port map (
            O => \N__3734\,
            I => char_42
        );

    \I__555\ : InMux
    port map (
            O => \N__3731\,
            I => \N__3728\
        );

    \I__554\ : LocalMux
    port map (
            O => \N__3728\,
            I => \tabla.n10\
        );

    \I__553\ : CascadeMux
    port map (
            O => \N__3725\,
            I => \tabla.n10_cascade_\
        );

    \I__552\ : CascadeMux
    port map (
            O => \N__3722\,
            I => \tabla.n1365_cascade_\
        );

    \I__551\ : CascadeMux
    port map (
            O => \N__3719\,
            I => \tabla.char_6_cascade_\
        );

    \I__550\ : CascadeMux
    port map (
            O => \N__3716\,
            I => \char_code_2_cascade_\
        );

    \I__549\ : InMux
    port map (
            O => \N__3713\,
            I => \N__3710\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__3710\,
            I => \generador.n1849\
        );

    \I__547\ : CascadeMux
    port map (
            O => \N__3707\,
            I => \n1949_cascade_\
        );

    \I__546\ : InMux
    port map (
            O => \N__3704\,
            I => \N__3701\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__3701\,
            I => \generador.n1958\
        );

    \I__544\ : InMux
    port map (
            O => \N__3698\,
            I => \N__3693\
        );

    \I__543\ : CascadeMux
    port map (
            O => \N__3697\,
            I => \N__3690\
        );

    \I__542\ : InMux
    port map (
            O => \N__3696\,
            I => \N__3687\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__3693\,
            I => \N__3683\
        );

    \I__540\ : InMux
    port map (
            O => \N__3690\,
            I => \N__3680\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__3687\,
            I => \N__3677\
        );

    \I__538\ : InMux
    port map (
            O => \N__3686\,
            I => \N__3674\
        );

    \I__537\ : Sp12to4
    port map (
            O => \N__3683\,
            I => \N__3666\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__3680\,
            I => \N__3666\
        );

    \I__535\ : Span4Mux_h
    port map (
            O => \N__3677\,
            I => \N__3661\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__3674\,
            I => \N__3661\
        );

    \I__533\ : InMux
    port map (
            O => \N__3673\,
            I => \N__3658\
        );

    \I__532\ : InMux
    port map (
            O => \N__3672\,
            I => \N__3653\
        );

    \I__531\ : InMux
    port map (
            O => \N__3671\,
            I => \N__3653\
        );

    \I__530\ : Odrv12
    port map (
            O => \N__3666\,
            I => linea_5
        );

    \I__529\ : Odrv4
    port map (
            O => \N__3661\,
            I => linea_5
        );

    \I__528\ : LocalMux
    port map (
            O => \N__3658\,
            I => linea_5
        );

    \I__527\ : LocalMux
    port map (
            O => \N__3653\,
            I => linea_5
        );

    \I__526\ : CascadeMux
    port map (
            O => \N__3644\,
            I => \N__3641\
        );

    \I__525\ : InMux
    port map (
            O => \N__3641\,
            I => \N__3638\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__3638\,
            I => \generador.n2000\
        );

    \I__523\ : CascadeMux
    port map (
            O => \N__3635\,
            I => \n1363_cascade_\
        );

    \I__522\ : CascadeMux
    port map (
            O => \N__3632\,
            I => \n1955_cascade_\
        );

    \I__521\ : InMux
    port map (
            O => \N__3629\,
            I => \N__3624\
        );

    \I__520\ : InMux
    port map (
            O => \N__3628\,
            I => \N__3615\
        );

    \I__519\ : InMux
    port map (
            O => \N__3627\,
            I => \N__3615\
        );

    \I__518\ : LocalMux
    port map (
            O => \N__3624\,
            I => \N__3612\
        );

    \I__517\ : InMux
    port map (
            O => \N__3623\,
            I => \N__3609\
        );

    \I__516\ : InMux
    port map (
            O => \N__3622\,
            I => \N__3602\
        );

    \I__515\ : InMux
    port map (
            O => \N__3621\,
            I => \N__3602\
        );

    \I__514\ : InMux
    port map (
            O => \N__3620\,
            I => \N__3602\
        );

    \I__513\ : LocalMux
    port map (
            O => \N__3615\,
            I => \N__3596\
        );

    \I__512\ : Span4Mux_v
    port map (
            O => \N__3612\,
            I => \N__3589\
        );

    \I__511\ : LocalMux
    port map (
            O => \N__3609\,
            I => \N__3589\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__3602\,
            I => \N__3589\
        );

    \I__509\ : InMux
    port map (
            O => \N__3601\,
            I => \N__3586\
        );

    \I__508\ : InMux
    port map (
            O => \N__3600\,
            I => \N__3581\
        );

    \I__507\ : InMux
    port map (
            O => \N__3599\,
            I => \N__3581\
        );

    \I__506\ : Odrv12
    port map (
            O => \N__3596\,
            I => linea_4
        );

    \I__505\ : Odrv4
    port map (
            O => \N__3589\,
            I => linea_4
        );

    \I__504\ : LocalMux
    port map (
            O => \N__3586\,
            I => linea_4
        );

    \I__503\ : LocalMux
    port map (
            O => \N__3581\,
            I => linea_4
        );

    \I__502\ : CascadeMux
    port map (
            O => \N__3572\,
            I => \generador.n1853_cascade_\
        );

    \I__501\ : InMux
    port map (
            O => \N__3569\,
            I => \N__3566\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__3566\,
            I => \generador.n1855\
        );

    \I__499\ : CascadeMux
    port map (
            O => \N__3563\,
            I => \tabla.char_57_cascade_\
        );

    \I__498\ : CascadeMux
    port map (
            O => \N__3560\,
            I => \n1399_cascade_\
        );

    \I__497\ : InMux
    port map (
            O => \N__3557\,
            I => \N__3546\
        );

    \I__496\ : InMux
    port map (
            O => \N__3556\,
            I => \N__3546\
        );

    \I__495\ : InMux
    port map (
            O => \N__3555\,
            I => \N__3546\
        );

    \I__494\ : InMux
    port map (
            O => \N__3554\,
            I => \N__3543\
        );

    \I__493\ : CascadeMux
    port map (
            O => \N__3553\,
            I => \N__3538\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__3546\,
            I => \N__3535\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__3543\,
            I => \N__3532\
        );

    \I__490\ : InMux
    port map (
            O => \N__3542\,
            I => \N__3529\
        );

    \I__489\ : InMux
    port map (
            O => \N__3541\,
            I => \N__3524\
        );

    \I__488\ : InMux
    port map (
            O => \N__3538\,
            I => \N__3524\
        );

    \I__487\ : Odrv4
    port map (
            O => \N__3535\,
            I => linea_6
        );

    \I__486\ : Odrv12
    port map (
            O => \N__3532\,
            I => linea_6
        );

    \I__485\ : LocalMux
    port map (
            O => \N__3529\,
            I => linea_6
        );

    \I__484\ : LocalMux
    port map (
            O => \N__3524\,
            I => linea_6
        );

    \I__483\ : CascadeMux
    port map (
            O => \N__3515\,
            I => \n32_cascade_\
        );

    \I__482\ : CascadeMux
    port map (
            O => \N__3512\,
            I => \generador.n1872_cascade_\
        );

    \I__481\ : InMux
    port map (
            O => \N__3509\,
            I => \N__3506\
        );

    \I__480\ : LocalMux
    port map (
            O => \N__3506\,
            I => \generador.n1961\
        );

    \I__479\ : InMux
    port map (
            O => \N__3503\,
            I => \N__3493\
        );

    \I__478\ : InMux
    port map (
            O => \N__3502\,
            I => \N__3493\
        );

    \I__477\ : InMux
    port map (
            O => \N__3501\,
            I => \N__3490\
        );

    \I__476\ : InMux
    port map (
            O => \N__3500\,
            I => \N__3485\
        );

    \I__475\ : InMux
    port map (
            O => \N__3499\,
            I => \N__3485\
        );

    \I__474\ : InMux
    port map (
            O => \N__3498\,
            I => \N__3482\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__3493\,
            I => n6
        );

    \I__472\ : LocalMux
    port map (
            O => \N__3490\,
            I => n6
        );

    \I__471\ : LocalMux
    port map (
            O => \N__3485\,
            I => n6
        );

    \I__470\ : LocalMux
    port map (
            O => \N__3482\,
            I => n6
        );

    \I__469\ : CascadeMux
    port map (
            O => \N__3473\,
            I => \N__3470\
        );

    \I__468\ : InMux
    port map (
            O => \N__3470\,
            I => \N__3464\
        );

    \I__467\ : InMux
    port map (
            O => \N__3469\,
            I => \N__3464\
        );

    \I__466\ : LocalMux
    port map (
            O => \N__3464\,
            I => \N__3455\
        );

    \I__465\ : InMux
    port map (
            O => \N__3463\,
            I => \N__3452\
        );

    \I__464\ : InMux
    port map (
            O => \N__3462\,
            I => \N__3447\
        );

    \I__463\ : InMux
    port map (
            O => \N__3461\,
            I => \N__3447\
        );

    \I__462\ : InMux
    port map (
            O => \N__3460\,
            I => \N__3440\
        );

    \I__461\ : InMux
    port map (
            O => \N__3459\,
            I => \N__3440\
        );

    \I__460\ : InMux
    port map (
            O => \N__3458\,
            I => \N__3440\
        );

    \I__459\ : Sp12to4
    port map (
            O => \N__3455\,
            I => \N__3432\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__3452\,
            I => \N__3432\
        );

    \I__457\ : LocalMux
    port map (
            O => \N__3447\,
            I => \N__3427\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__3440\,
            I => \N__3427\
        );

    \I__455\ : InMux
    port map (
            O => \N__3439\,
            I => \N__3424\
        );

    \I__454\ : InMux
    port map (
            O => \N__3438\,
            I => \N__3421\
        );

    \I__453\ : InMux
    port map (
            O => \N__3437\,
            I => \N__3418\
        );

    \I__452\ : Odrv12
    port map (
            O => \N__3432\,
            I => linea_7
        );

    \I__451\ : Odrv4
    port map (
            O => \N__3427\,
            I => linea_7
        );

    \I__450\ : LocalMux
    port map (
            O => \N__3424\,
            I => linea_7
        );

    \I__449\ : LocalMux
    port map (
            O => \N__3421\,
            I => linea_7
        );

    \I__448\ : LocalMux
    port map (
            O => \N__3418\,
            I => linea_7
        );

    \I__447\ : InMux
    port map (
            O => \N__3407\,
            I => \N__3400\
        );

    \I__446\ : InMux
    port map (
            O => \N__3406\,
            I => \N__3400\
        );

    \I__445\ : CascadeMux
    port map (
            O => \N__3405\,
            I => \N__3395\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__3400\,
            I => \N__3390\
        );

    \I__443\ : InMux
    port map (
            O => \N__3399\,
            I => \N__3387\
        );

    \I__442\ : InMux
    port map (
            O => \N__3398\,
            I => \N__3384\
        );

    \I__441\ : InMux
    port map (
            O => \N__3395\,
            I => \N__3379\
        );

    \I__440\ : InMux
    port map (
            O => \N__3394\,
            I => \N__3379\
        );

    \I__439\ : InMux
    port map (
            O => \N__3393\,
            I => \N__3373\
        );

    \I__438\ : Span4Mux_h
    port map (
            O => \N__3390\,
            I => \N__3364\
        );

    \I__437\ : LocalMux
    port map (
            O => \N__3387\,
            I => \N__3364\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__3384\,
            I => \N__3364\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__3379\,
            I => \N__3364\
        );

    \I__434\ : InMux
    port map (
            O => \N__3378\,
            I => \N__3361\
        );

    \I__433\ : InMux
    port map (
            O => \N__3377\,
            I => \N__3356\
        );

    \I__432\ : InMux
    port map (
            O => \N__3376\,
            I => \N__3356\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__3373\,
            I => linea_8
        );

    \I__430\ : Odrv4
    port map (
            O => \N__3364\,
            I => linea_8
        );

    \I__429\ : LocalMux
    port map (
            O => \N__3361\,
            I => linea_8
        );

    \I__428\ : LocalMux
    port map (
            O => \N__3356\,
            I => linea_8
        );

    \I__427\ : CascadeMux
    port map (
            O => \N__3347\,
            I => \n1946_cascade_\
        );

    \I__426\ : InMux
    port map (
            O => \N__3344\,
            I => \sincronismo.n1569\
        );

    \I__425\ : InMux
    port map (
            O => \N__3341\,
            I => \bfn_6_12_0_\
        );

    \I__424\ : InMux
    port map (
            O => \N__3338\,
            I => \sincronismo.n1571\
        );

    \I__423\ : InMux
    port map (
            O => \N__3335\,
            I => \N__3331\
        );

    \I__422\ : CascadeMux
    port map (
            O => \N__3334\,
            I => \N__3327\
        );

    \I__421\ : LocalMux
    port map (
            O => \N__3331\,
            I => \N__3323\
        );

    \I__420\ : InMux
    port map (
            O => \N__3330\,
            I => \N__3320\
        );

    \I__419\ : InMux
    port map (
            O => \N__3327\,
            I => \N__3315\
        );

    \I__418\ : InMux
    port map (
            O => \N__3326\,
            I => \N__3315\
        );

    \I__417\ : Odrv4
    port map (
            O => \N__3323\,
            I => linea_9
        );

    \I__416\ : LocalMux
    port map (
            O => \N__3320\,
            I => linea_9
        );

    \I__415\ : LocalMux
    port map (
            O => \N__3315\,
            I => linea_9
        );

    \I__414\ : ClkMux
    port map (
            O => \N__3308\,
            I => \N__3296\
        );

    \I__413\ : ClkMux
    port map (
            O => \N__3307\,
            I => \N__3296\
        );

    \I__412\ : ClkMux
    port map (
            O => \N__3306\,
            I => \N__3296\
        );

    \I__411\ : ClkMux
    port map (
            O => \N__3305\,
            I => \N__3296\
        );

    \I__410\ : GlobalMux
    port map (
            O => \N__3296\,
            I => p_clk
        );

    \I__409\ : CEMux
    port map (
            O => \N__3293\,
            I => \N__3290\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__3290\,
            I => \N__3285\
        );

    \I__407\ : SRMux
    port map (
            O => \N__3289\,
            I => \N__3281\
        );

    \I__406\ : SRMux
    port map (
            O => \N__3288\,
            I => \N__3278\
        );

    \I__405\ : Span4Mux_v
    port map (
            O => \N__3285\,
            I => \N__3275\
        );

    \I__404\ : CEMux
    port map (
            O => \N__3284\,
            I => \N__3272\
        );

    \I__403\ : LocalMux
    port map (
            O => \N__3281\,
            I => \N__3269\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__3278\,
            I => \N__3266\
        );

    \I__401\ : Span4Mux_v
    port map (
            O => \N__3275\,
            I => \N__3261\
        );

    \I__400\ : LocalMux
    port map (
            O => \N__3272\,
            I => \N__3261\
        );

    \I__399\ : Span4Mux_v
    port map (
            O => \N__3269\,
            I => \N__3258\
        );

    \I__398\ : Span4Mux_h
    port map (
            O => \N__3266\,
            I => \N__3255\
        );

    \I__397\ : Odrv4
    port map (
            O => \N__3261\,
            I => \sincronismo.n1006\
        );

    \I__396\ : Odrv4
    port map (
            O => \N__3258\,
            I => \sincronismo.n1006\
        );

    \I__395\ : Odrv4
    port map (
            O => \N__3255\,
            I => \sincronismo.n1006\
        );

    \I__394\ : SRMux
    port map (
            O => \N__3248\,
            I => \N__3245\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__3245\,
            I => \N__3241\
        );

    \I__392\ : SRMux
    port map (
            O => \N__3244\,
            I => \N__3238\
        );

    \I__391\ : Span4Mux_h
    port map (
            O => \N__3241\,
            I => \N__3233\
        );

    \I__390\ : LocalMux
    port map (
            O => \N__3238\,
            I => \N__3233\
        );

    \I__389\ : Odrv4
    port map (
            O => \N__3233\,
            I => \sincronismo.n1033\
        );

    \I__388\ : CascadeMux
    port map (
            O => \N__3230\,
            I => \N__3227\
        );

    \I__387\ : InMux
    port map (
            O => \N__3227\,
            I => \N__3224\
        );

    \I__386\ : LocalMux
    port map (
            O => \N__3224\,
            I => \sincronismo.n1884\
        );

    \I__385\ : CascadeMux
    port map (
            O => \N__3221\,
            I => \sincronismo.n1932_cascade_\
        );

    \I__384\ : CascadeMux
    port map (
            O => \N__3218\,
            I => \N__3215\
        );

    \I__383\ : InMux
    port map (
            O => \N__3215\,
            I => \N__3212\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__3212\,
            I => n14_adj_135
        );

    \I__381\ : InMux
    port map (
            O => \N__3209\,
            I => \N__3199\
        );

    \I__380\ : InMux
    port map (
            O => \N__3208\,
            I => \N__3199\
        );

    \I__379\ : InMux
    port map (
            O => \N__3207\,
            I => \N__3199\
        );

    \I__378\ : InMux
    port map (
            O => \N__3206\,
            I => \N__3196\
        );

    \I__377\ : LocalMux
    port map (
            O => \N__3199\,
            I => n1928
        );

    \I__376\ : LocalMux
    port map (
            O => \N__3196\,
            I => n1928
        );

    \I__375\ : CascadeMux
    port map (
            O => \N__3191\,
            I => \n1928_cascade_\
        );

    \I__374\ : InMux
    port map (
            O => \N__3188\,
            I => \N__3182\
        );

    \I__373\ : InMux
    port map (
            O => \N__3187\,
            I => \N__3182\
        );

    \I__372\ : LocalMux
    port map (
            O => \N__3182\,
            I => linea_z_1
        );

    \I__371\ : InMux
    port map (
            O => \N__3179\,
            I => \N__3175\
        );

    \I__370\ : InMux
    port map (
            O => \N__3178\,
            I => \N__3172\
        );

    \I__369\ : LocalMux
    port map (
            O => \N__3175\,
            I => \N__3167\
        );

    \I__368\ : LocalMux
    port map (
            O => \N__3172\,
            I => \N__3167\
        );

    \I__367\ : Odrv4
    port map (
            O => \N__3167\,
            I => \sincronismo.linea_0\
        );

    \I__366\ : InMux
    port map (
            O => \N__3164\,
            I => \bfn_6_11_0_\
        );

    \I__365\ : CascadeMux
    port map (
            O => \N__3161\,
            I => \N__3157\
        );

    \I__364\ : InMux
    port map (
            O => \N__3160\,
            I => \N__3153\
        );

    \I__363\ : InMux
    port map (
            O => \N__3157\,
            I => \N__3148\
        );

    \I__362\ : InMux
    port map (
            O => \N__3156\,
            I => \N__3148\
        );

    \I__361\ : LocalMux
    port map (
            O => \N__3153\,
            I => \sincronismo.linea_1\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__3148\,
            I => \sincronismo.linea_1\
        );

    \I__359\ : InMux
    port map (
            O => \N__3143\,
            I => \sincronismo.n1563\
        );

    \I__358\ : InMux
    port map (
            O => \N__3140\,
            I => \N__3135\
        );

    \I__357\ : InMux
    port map (
            O => \N__3139\,
            I => \N__3132\
        );

    \I__356\ : InMux
    port map (
            O => \N__3138\,
            I => \N__3129\
        );

    \I__355\ : LocalMux
    port map (
            O => \N__3135\,
            I => \sincronismo.linea_2\
        );

    \I__354\ : LocalMux
    port map (
            O => \N__3132\,
            I => \sincronismo.linea_2\
        );

    \I__353\ : LocalMux
    port map (
            O => \N__3129\,
            I => \sincronismo.linea_2\
        );

    \I__352\ : InMux
    port map (
            O => \N__3122\,
            I => \sincronismo.n1564\
        );

    \I__351\ : InMux
    port map (
            O => \N__3119\,
            I => \N__3114\
        );

    \I__350\ : InMux
    port map (
            O => \N__3118\,
            I => \N__3109\
        );

    \I__349\ : InMux
    port map (
            O => \N__3117\,
            I => \N__3109\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__3114\,
            I => \sincronismo.linea_3\
        );

    \I__347\ : LocalMux
    port map (
            O => \N__3109\,
            I => \sincronismo.linea_3\
        );

    \I__346\ : InMux
    port map (
            O => \N__3104\,
            I => \sincronismo.n1565\
        );

    \I__345\ : InMux
    port map (
            O => \N__3101\,
            I => \sincronismo.n1566\
        );

    \I__344\ : InMux
    port map (
            O => \N__3098\,
            I => \sincronismo.n1567\
        );

    \I__343\ : InMux
    port map (
            O => \N__3095\,
            I => \sincronismo.n1568\
        );

    \I__342\ : InMux
    port map (
            O => \N__3092\,
            I => \N__3089\
        );

    \I__341\ : LocalMux
    port map (
            O => \N__3089\,
            I => \salida.n1886\
        );

    \I__340\ : CascadeMux
    port map (
            O => \N__3086\,
            I => \generador.n2003_cascade_\
        );

    \I__339\ : CascadeMux
    port map (
            O => \N__3083\,
            I => \generador.px_visible_N_105_cascade_\
        );

    \I__338\ : IoInMux
    port map (
            O => \N__3080\,
            I => \N__3077\
        );

    \I__337\ : LocalMux
    port map (
            O => \N__3077\,
            I => \N__3074\
        );

    \I__336\ : Span4Mux_s1_h
    port map (
            O => \N__3074\,
            I => \N__3071\
        );

    \I__335\ : Sp12to4
    port map (
            O => \N__3071\,
            I => \N__3068\
        );

    \I__334\ : Span12Mux_v
    port map (
            O => \N__3068\,
            I => \N__3065\
        );

    \I__333\ : Odrv12
    port map (
            O => \N__3065\,
            I => pixel_c
        );

    \I__332\ : InMux
    port map (
            O => \N__3062\,
            I => \N__3059\
        );

    \I__331\ : LocalMux
    port map (
            O => \N__3059\,
            I => \generador.n1856\
        );

    \I__330\ : InMux
    port map (
            O => \N__3056\,
            I => \N__3053\
        );

    \I__329\ : LocalMux
    port map (
            O => \N__3053\,
            I => \generador.n1843\
        );

    \I__328\ : CascadeMux
    port map (
            O => \N__3050\,
            I => \N__3046\
        );

    \I__327\ : InMux
    port map (
            O => \N__3049\,
            I => \N__3038\
        );

    \I__326\ : InMux
    port map (
            O => \N__3046\,
            I => \N__3038\
        );

    \I__325\ : InMux
    port map (
            O => \N__3045\,
            I => \N__3038\
        );

    \I__324\ : LocalMux
    port map (
            O => \N__3038\,
            I => n517
        );

    \I__323\ : CascadeMux
    port map (
            O => \N__3035\,
            I => \n1001_cascade_\
        );

    \I__322\ : InMux
    port map (
            O => \N__3032\,
            I => \N__3027\
        );

    \I__321\ : InMux
    port map (
            O => \N__3031\,
            I => \N__3022\
        );

    \I__320\ : InMux
    port map (
            O => \N__3030\,
            I => \N__3022\
        );

    \I__319\ : LocalMux
    port map (
            O => \N__3027\,
            I => n1167
        );

    \I__318\ : LocalMux
    port map (
            O => \N__3022\,
            I => n1167
        );

    \I__317\ : InMux
    port map (
            O => \N__3017\,
            I => \N__3014\
        );

    \I__316\ : LocalMux
    port map (
            O => \N__3014\,
            I => \generador.n6\
        );

    \I__315\ : CascadeMux
    port map (
            O => \N__3011\,
            I => \n14_adj_131_cascade_\
        );

    \I__314\ : InMux
    port map (
            O => \N__3008\,
            I => \N__3005\
        );

    \I__313\ : LocalMux
    port map (
            O => \N__3005\,
            I => \sincronismo.n1839\
        );

    \I__312\ : CascadeMux
    port map (
            O => \N__3002\,
            I => \sincronismo.n1006_cascade_\
        );

    \I__311\ : InMux
    port map (
            O => \N__2999\,
            I => \N__2996\
        );

    \I__310\ : LocalMux
    port map (
            O => \N__2996\,
            I => \sincronismo.n10\
        );

    \I__309\ : InMux
    port map (
            O => \N__2993\,
            I => \N__2989\
        );

    \I__308\ : InMux
    port map (
            O => \N__2992\,
            I => \N__2986\
        );

    \I__307\ : LocalMux
    port map (
            O => \N__2989\,
            I => \sincronismo.n1823\
        );

    \I__306\ : LocalMux
    port map (
            O => \N__2986\,
            I => \sincronismo.n1823\
        );

    \I__305\ : InMux
    port map (
            O => \N__2981\,
            I => \N__2978\
        );

    \I__304\ : LocalMux
    port map (
            O => \N__2978\,
            I => \sincronismo.n1401\
        );

    \I__303\ : InMux
    port map (
            O => \N__2975\,
            I => \N__2969\
        );

    \I__302\ : InMux
    port map (
            O => \N__2974\,
            I => \N__2969\
        );

    \I__301\ : LocalMux
    port map (
            O => \N__2969\,
            I => \sincronismo.n980\
        );

    \I__300\ : IoInMux
    port map (
            O => \N__2966\,
            I => \N__2963\
        );

    \I__299\ : LocalMux
    port map (
            O => \N__2963\,
            I => \N__2960\
        );

    \I__298\ : IoSpan4Mux
    port map (
            O => \N__2960\,
            I => \N__2957\
        );

    \I__297\ : Span4Mux_s1_h
    port map (
            O => \N__2957\,
            I => \N__2954\
        );

    \I__296\ : Sp12to4
    port map (
            O => \N__2954\,
            I => \N__2951\
        );

    \I__295\ : Span12Mux_s8_h
    port map (
            O => \N__2951\,
            I => \N__2948\
        );

    \I__294\ : Odrv12
    port map (
            O => \N__2948\,
            I => \vsync_N_90\
        );

    \I__293\ : CascadeMux
    port map (
            O => \N__2945\,
            I => \n15_adj_136_cascade_\
        );

    \I__292\ : CascadeMux
    port map (
            O => \N__2942\,
            I => \sincronismo.n1890_cascade_\
        );

    \I__291\ : InMux
    port map (
            O => \N__2939\,
            I => \N__2936\
        );

    \I__290\ : LocalMux
    port map (
            O => \N__2936\,
            I => \sincronismo.n51\
        );

    \I__289\ : CascadeMux
    port map (
            O => \N__2933\,
            I => \sincronismo.n1889_cascade_\
        );

    \I__288\ : InMux
    port map (
            O => \N__2930\,
            I => \N__2927\
        );

    \I__287\ : LocalMux
    port map (
            O => \N__2927\,
            I => \sincronismo.n1193\
        );

    \I__286\ : IoInMux
    port map (
            O => \N__2924\,
            I => \N__2921\
        );

    \I__285\ : LocalMux
    port map (
            O => \N__2921\,
            I => \N__2918\
        );

    \I__284\ : IoSpan4Mux
    port map (
            O => \N__2918\,
            I => \N__2915\
        );

    \I__283\ : Span4Mux_s2_h
    port map (
            O => \N__2915\,
            I => \N__2912\
        );

    \I__282\ : Span4Mux_h
    port map (
            O => \N__2912\,
            I => \N__2909\
        );

    \I__281\ : Odrv4
    port map (
            O => \N__2909\,
            I => h_sync_c
        );

    \I__280\ : CascadeMux
    port map (
            O => \N__2906\,
            I => \sincronismo.n1383_cascade_\
        );

    \I__279\ : CascadeMux
    port map (
            O => \N__2903\,
            I => \sincronismo.n6_cascade_\
        );

    \I__278\ : CascadeMux
    port map (
            O => \N__2900\,
            I => \N__2896\
        );

    \I__277\ : InMux
    port map (
            O => \N__2899\,
            I => \N__2893\
        );

    \I__276\ : InMux
    port map (
            O => \N__2896\,
            I => \N__2889\
        );

    \I__275\ : LocalMux
    port map (
            O => \N__2893\,
            I => \N__2886\
        );

    \I__274\ : InMux
    port map (
            O => \N__2892\,
            I => \N__2883\
        );

    \I__273\ : LocalMux
    port map (
            O => \N__2889\,
            I => \N__2880\
        );

    \I__272\ : Odrv12
    port map (
            O => \N__2886\,
            I => columna_3
        );

    \I__271\ : LocalMux
    port map (
            O => \N__2883\,
            I => columna_3
        );

    \I__270\ : Odrv4
    port map (
            O => \N__2880\,
            I => columna_3
        );

    \I__269\ : InMux
    port map (
            O => \N__2873\,
            I => \N__2870\
        );

    \I__268\ : LocalMux
    port map (
            O => \N__2870\,
            I => \N__2867\
        );

    \I__267\ : Span4Mux_h
    port map (
            O => \N__2867\,
            I => \N__2864\
        );

    \I__266\ : Odrv4
    port map (
            O => \N__2864\,
            I => n1809
        );

    \I__265\ : InMux
    port map (
            O => \N__2861\,
            I => \sincronismo.n1573\
        );

    \I__264\ : InMux
    port map (
            O => \N__2858\,
            I => \sincronismo.n1574\
        );

    \I__263\ : InMux
    port map (
            O => \N__2855\,
            I => \sincronismo.n1575\
        );

    \I__262\ : InMux
    port map (
            O => \N__2852\,
            I => \sincronismo.n1576\
        );

    \I__261\ : InMux
    port map (
            O => \N__2849\,
            I => \sincronismo.n1577\
        );

    \I__260\ : InMux
    port map (
            O => \N__2846\,
            I => \sincronismo.n1578\
        );

    \I__259\ : InMux
    port map (
            O => \N__2843\,
            I => \bfn_3_13_0_\
        );

    \I__258\ : InMux
    port map (
            O => \N__2840\,
            I => \sincronismo.n1580\
        );

    \I__257\ : InMux
    port map (
            O => \N__2837\,
            I => \N__2833\
        );

    \I__256\ : CascadeMux
    port map (
            O => \N__2836\,
            I => \N__2829\
        );

    \I__255\ : LocalMux
    port map (
            O => \N__2833\,
            I => \N__2826\
        );

    \I__254\ : InMux
    port map (
            O => \N__2832\,
            I => \N__2823\
        );

    \I__253\ : InMux
    port map (
            O => \N__2829\,
            I => \N__2820\
        );

    \I__252\ : Odrv4
    port map (
            O => \N__2826\,
            I => \sincronismo.columna_1\
        );

    \I__251\ : LocalMux
    port map (
            O => \N__2823\,
            I => \sincronismo.columna_1\
        );

    \I__250\ : LocalMux
    port map (
            O => \N__2820\,
            I => \sincronismo.columna_1\
        );

    \I__249\ : CascadeMux
    port map (
            O => \N__2813\,
            I => \N__2810\
        );

    \I__248\ : InMux
    port map (
            O => \N__2810\,
            I => \N__2807\
        );

    \I__247\ : LocalMux
    port map (
            O => \N__2807\,
            I => \N__2802\
        );

    \I__246\ : InMux
    port map (
            O => \N__2806\,
            I => \N__2799\
        );

    \I__245\ : InMux
    port map (
            O => \N__2805\,
            I => \N__2796\
        );

    \I__244\ : Odrv12
    port map (
            O => \N__2802\,
            I => \sincronismo.columna_0\
        );

    \I__243\ : LocalMux
    port map (
            O => \N__2799\,
            I => \sincronismo.columna_0\
        );

    \I__242\ : LocalMux
    port map (
            O => \N__2796\,
            I => \sincronismo.columna_0\
        );

    \I__241\ : InMux
    port map (
            O => \N__2789\,
            I => \N__2786\
        );

    \I__240\ : LocalMux
    port map (
            O => \N__2786\,
            I => \N__2781\
        );

    \I__239\ : InMux
    port map (
            O => \N__2785\,
            I => \N__2778\
        );

    \I__238\ : InMux
    port map (
            O => \N__2784\,
            I => \N__2775\
        );

    \I__237\ : Odrv4
    port map (
            O => \N__2781\,
            I => \sincronismo.columna_2\
        );

    \I__236\ : LocalMux
    port map (
            O => \N__2778\,
            I => \sincronismo.columna_2\
        );

    \I__235\ : LocalMux
    port map (
            O => \N__2775\,
            I => \sincronismo.columna_2\
        );

    \I__234\ : InMux
    port map (
            O => \N__2768\,
            I => \bfn_3_12_0_\
        );

    \I__233\ : InMux
    port map (
            O => \N__2765\,
            I => \sincronismo.n1572\
        );

    \IN_MUX_bfv_6_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_11_0_\
        );

    \IN_MUX_bfv_6_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sincronismo.n1570\,
            carryinitout => \bfn_6_12_0_\
        );

    \IN_MUX_bfv_3_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_3_12_0_\
        );

    \IN_MUX_bfv_3_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \sincronismo.n1579\,
            carryinitout => \bfn_3_13_0_\
        );

    \IN_MUX_bfv_12_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_11_0_\
        );

    \IN_MUX_bfv_12_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n1539,
            carryinitout => \bfn_12_12_0_\
        );

    \IN_MUX_bfv_12_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n1547,
            carryinitout => \bfn_12_13_0_\
        );

    \IN_MUX_bfv_12_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => n1555,
            carryinitout => \bfn_12_14_0_\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \sincronismo.i2_3_lut_adj_6_LC_3_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010000000"
        )
    port map (
            in0 => \N__2805\,
            in1 => \N__2784\,
            in2 => \N__2836\,
            in3 => \_gnd_net_\,
            lcout => n1809,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.Q_46__i0_LC_3_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2806\,
            in2 => \_gnd_net_\,
            in3 => \N__2768\,
            lcout => \sincronismo.columna_0\,
            ltout => OPEN,
            carryin => \bfn_3_12_0_\,
            carryout => \sincronismo.n1572\,
            clk => \N__3307\,
            ce => 'H',
            sr => \N__3288\
        );

    \sincronismo.Q_46__i1_LC_3_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2832\,
            in2 => \_gnd_net_\,
            in3 => \N__2765\,
            lcout => \sincronismo.columna_1\,
            ltout => OPEN,
            carryin => \sincronismo.n1572\,
            carryout => \sincronismo.n1573\,
            clk => \N__3307\,
            ce => 'H',
            sr => \N__3288\
        );

    \sincronismo.Q_46__i2_LC_3_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2785\,
            in2 => \_gnd_net_\,
            in3 => \N__2861\,
            lcout => \sincronismo.columna_2\,
            ltout => OPEN,
            carryin => \sincronismo.n1573\,
            carryout => \sincronismo.n1574\,
            clk => \N__3307\,
            ce => 'H',
            sr => \N__3288\
        );

    \sincronismo.Q_46__i3_LC_3_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__2892\,
            in2 => \_gnd_net_\,
            in3 => \N__2858\,
            lcout => columna_3,
            ltout => OPEN,
            carryin => \sincronismo.n1574\,
            carryout => \sincronismo.n1575\,
            clk => \N__3307\,
            ce => 'H',
            sr => \N__3288\
        );

    \sincronismo.Q_46__i4_LC_3_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4899\,
            in2 => \_gnd_net_\,
            in3 => \N__2855\,
            lcout => columna_4,
            ltout => OPEN,
            carryin => \sincronismo.n1575\,
            carryout => \sincronismo.n1576\,
            clk => \N__3307\,
            ce => 'H',
            sr => \N__3288\
        );

    \sincronismo.Q_46__i5_LC_3_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5933\,
            in2 => \_gnd_net_\,
            in3 => \N__2852\,
            lcout => columna_5,
            ltout => OPEN,
            carryin => \sincronismo.n1576\,
            carryout => \sincronismo.n1577\,
            clk => \N__3307\,
            ce => 'H',
            sr => \N__3288\
        );

    \sincronismo.Q_46__i6_LC_3_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4469\,
            in2 => \_gnd_net_\,
            in3 => \N__2849\,
            lcout => columna_6,
            ltout => OPEN,
            carryin => \sincronismo.n1577\,
            carryout => \sincronismo.n1578\,
            clk => \N__3307\,
            ce => 'H',
            sr => \N__3288\
        );

    \sincronismo.Q_46__i7_LC_3_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3804\,
            in2 => \_gnd_net_\,
            in3 => \N__2846\,
            lcout => columna_7,
            ltout => OPEN,
            carryin => \sincronismo.n1578\,
            carryout => \sincronismo.n1579\,
            clk => \N__3307\,
            ce => 'H',
            sr => \N__3288\
        );

    \sincronismo.Q_46__i8_LC_3_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4757\,
            in2 => \_gnd_net_\,
            in3 => \N__2843\,
            lcout => columna_8,
            ltout => OPEN,
            carryin => \bfn_3_13_0_\,
            carryout => \sincronismo.n1580\,
            clk => \N__3308\,
            ce => 'H',
            sr => \N__3289\
        );

    \sincronismo.Q_46__i9_LC_3_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4643\,
            in2 => \_gnd_net_\,
            in3 => \N__2840\,
            lcout => columna_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3308\,
            ce => 'H',
            sr => \N__3289\
        );

    \sincronismo.i1446_2_lut_4_lut_LC_3_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__2837\,
            in1 => \N__2899\,
            in2 => \N__2813\,
            in3 => \N__2789\,
            lcout => OPEN,
            ltout => \sincronismo.n1889_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i803_4_lut_LC_3_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000010001"
        )
    port map (
            in0 => \N__5971\,
            in1 => \N__4938\,
            in2 => \N__2933\,
            in3 => \N__4476\,
            lcout => \sincronismo.n1193\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i2_4_lut_LC_3_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__2930\,
            in1 => \N__4677\,
            in2 => \N__4820\,
            in3 => \N__3815\,
            lcout => h_sync_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i989_4_lut_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011001100"
        )
    port map (
            in0 => \N__2992\,
            in1 => \N__3672\,
            in2 => \N__3161\,
            in3 => \N__3600\,
            lcout => OPEN,
            ltout => \sincronismo.n1383_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i1003_4_lut_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__3541\,
            in1 => \N__3439\,
            in2 => \N__2906\,
            in3 => \N__3377\,
            lcout => \sincronismo.n1401\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i1_2_lut_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__3118\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3140\,
            lcout => \sincronismo.n1823\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i1_2_lut_4_lut_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3437\,
            in1 => \N__3376\,
            in2 => \N__3553\,
            in3 => \N__3156\,
            lcout => OPEN,
            ltout => \sincronismo.n6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i4_4_lut_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3178\,
            in1 => \N__3671\,
            in2 => \N__2903\,
            in3 => \N__3599\,
            lcout => \sincronismo.n980\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i1376_2_lut_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3117\,
            in2 => \_gnd_net_\,
            in3 => \N__3138\,
            lcout => \sincronismo.n1839\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generador.i6_4_lut_4_lut_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__4806\,
            in1 => \N__5950\,
            in2 => \N__2900\,
            in3 => \N__2873\,
            lcout => OPEN,
            ltout => \n14_adj_131_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i7_4_lut_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__4696\,
            in1 => \N__4468\,
            in2 => \N__3011\,
            in3 => \N__2999\,
            lcout => \sincronismo.n1006\,
            ltout => \sincronismo.n1006_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i641_4_lut_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__3326\,
            in1 => \N__3008\,
            in2 => \N__3002\,
            in3 => \N__2974\,
            lcout => \sincronismo.n1033\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i2_2_lut_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3803\,
            in2 => \_gnd_net_\,
            in3 => \N__4912\,
            lcout => \sincronismo.n10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i1475_4_lut_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111111011111"
        )
    port map (
            in0 => \N__2993\,
            in1 => \N__2981\,
            in2 => \N__3334\,
            in3 => \N__2975\,
            lcout => \vsync_N_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \salida.n_zona_4__I_0_Mux_1_i15_4_lut_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010111011"
        )
    port map (
            in0 => \N__3092\,
            in1 => \N__3207\,
            in2 => \N__3218\,
            in3 => \N__4807\,
            lcout => OPEN,
            ltout => \n15_adj_136_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i1_4_lut_adj_5_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111111100"
        )
    port map (
            in0 => \N__3209\,
            in1 => \N__3031\,
            in2 => \N__2945\,
            in3 => \N__4699\,
            lcout => char_code_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i1460_2_lut_3_lut_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011011101"
        )
    port map (
            in0 => \N__3503\,
            in1 => \N__3393\,
            in2 => \_gnd_net_\,
            in3 => \N__3462\,
            lcout => OPEN,
            ltout => \sincronismo.n1890_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i1_4_lut_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111010001"
        )
    port map (
            in0 => \N__3208\,
            in1 => \N__2939\,
            in2 => \N__2942\,
            in3 => \N__3030\,
            lcout => char_code_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i1_3_lut_adj_9_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010101010"
        )
    port map (
            in0 => \N__4698\,
            in1 => \_gnd_net_\,
            in2 => \N__3832\,
            in3 => \N__4809\,
            lcout => \sincronismo.n51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \salida.i1453_2_lut_3_lut_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100100000000"
        )
    port map (
            in0 => \N__3461\,
            in1 => \N__3502\,
            in2 => \_gnd_net_\,
            in3 => \N__3822\,
            lcout => \salida.n1886\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i1_3_lut_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010001000"
        )
    port map (
            in0 => \N__4808\,
            in1 => \N__4697\,
            in2 => \_gnd_net_\,
            in3 => \N__3823\,
            lcout => n1167,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \posicion.i122_2_lut_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__3623\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3696\,
            lcout => n517,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generador.n2000_bdd_4_lut_4_lut_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101011010000"
        )
    port map (
            in0 => \N__3188\,
            in1 => \N__3983\,
            in2 => \N__3644\,
            in3 => \N__4079\,
            lcout => OPEN,
            ltout => \generador.n2003_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generador.i104914_i1_4_lut_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010111000"
        )
    port map (
            in0 => \N__3062\,
            in1 => \N__3045\,
            in2 => \N__3086\,
            in3 => \N__3555\,
            lcout => OPEN,
            ltout => \generador.px_visible_N_105_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generador.i4_4_lut_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__3056\,
            in1 => \N__3017\,
            in2 => \N__3083\,
            in3 => \N__3335\,
            lcout => pixel_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generador.i1393_3_lut_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__3509\,
            in1 => \N__3187\,
            in2 => \_gnd_net_\,
            in3 => \N__3569\,
            lcout => \generador.n1856\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generador.i1380_3_lut_4_lut_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000000000"
        )
    port map (
            in0 => \N__3556\,
            in1 => \N__3469\,
            in2 => \N__3050\,
            in3 => \N__3406\,
            lcout => \generador.n1843\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i2_3_lut_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111010"
        )
    port map (
            in0 => \N__3407\,
            in1 => \_gnd_net_\,
            in2 => \N__3473\,
            in3 => \N__3557\,
            lcout => OPEN,
            ltout => \n1001_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generador.i1_3_lut_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111010"
        )
    port map (
            in0 => \N__3049\,
            in1 => \_gnd_net_\,
            in2 => \N__3035\,
            in3 => \N__3032\,
            lcout => \generador.n6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \posicion.i120_2_lut_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3698\,
            in2 => \_gnd_net_\,
            in3 => \N__3629\,
            lcout => linea_z_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.Q_47__i0_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3179\,
            in2 => \_gnd_net_\,
            in3 => \N__3164\,
            lcout => \sincronismo.linea_0\,
            ltout => OPEN,
            carryin => \bfn_6_11_0_\,
            carryout => \sincronismo.n1563\,
            clk => \N__3305\,
            ce => \N__3293\,
            sr => \N__3248\
        );

    \sincronismo.Q_47__i1_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3160\,
            in2 => \_gnd_net_\,
            in3 => \N__3143\,
            lcout => \sincronismo.linea_1\,
            ltout => OPEN,
            carryin => \sincronismo.n1563\,
            carryout => \sincronismo.n1564\,
            clk => \N__3305\,
            ce => \N__3293\,
            sr => \N__3248\
        );

    \sincronismo.Q_47__i2_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3139\,
            in2 => \_gnd_net_\,
            in3 => \N__3122\,
            lcout => \sincronismo.linea_2\,
            ltout => OPEN,
            carryin => \sincronismo.n1564\,
            carryout => \sincronismo.n1565\,
            clk => \N__3305\,
            ce => \N__3293\,
            sr => \N__3248\
        );

    \sincronismo.Q_47__i3_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3119\,
            in2 => \_gnd_net_\,
            in3 => \N__3104\,
            lcout => \sincronismo.linea_3\,
            ltout => OPEN,
            carryin => \sincronismo.n1565\,
            carryout => \sincronismo.n1566\,
            clk => \N__3305\,
            ce => \N__3293\,
            sr => \N__3248\
        );

    \sincronismo.Q_47__i4_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3601\,
            in2 => \_gnd_net_\,
            in3 => \N__3101\,
            lcout => linea_4,
            ltout => OPEN,
            carryin => \sincronismo.n1566\,
            carryout => \sincronismo.n1567\,
            clk => \N__3305\,
            ce => \N__3293\,
            sr => \N__3248\
        );

    \sincronismo.Q_47__i5_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3673\,
            in2 => \_gnd_net_\,
            in3 => \N__3098\,
            lcout => linea_5,
            ltout => OPEN,
            carryin => \sincronismo.n1567\,
            carryout => \sincronismo.n1568\,
            clk => \N__3305\,
            ce => \N__3293\,
            sr => \N__3248\
        );

    \sincronismo.Q_47__i6_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3542\,
            in2 => \_gnd_net_\,
            in3 => \N__3095\,
            lcout => linea_6,
            ltout => OPEN,
            carryin => \sincronismo.n1568\,
            carryout => \sincronismo.n1569\,
            clk => \N__3305\,
            ce => \N__3293\,
            sr => \N__3248\
        );

    \sincronismo.Q_47__i7_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3438\,
            in2 => \_gnd_net_\,
            in3 => \N__3344\,
            lcout => linea_7,
            ltout => OPEN,
            carryin => \sincronismo.n1569\,
            carryout => \sincronismo.n1570\,
            clk => \N__3305\,
            ce => \N__3293\,
            sr => \N__3248\
        );

    \sincronismo.Q_47__i8_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3378\,
            in2 => \_gnd_net_\,
            in3 => \N__3341\,
            lcout => linea_8,
            ltout => OPEN,
            carryin => \bfn_6_12_0_\,
            carryout => \sincronismo.n1571\,
            clk => \N__3306\,
            ce => \N__3284\,
            sr => \N__3244\
        );

    \sincronismo.Q_47__i9_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3330\,
            in2 => \_gnd_net_\,
            in3 => \N__3338\,
            lcout => linea_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__3306\,
            ce => \N__3284\,
            sr => \N__3244\
        );

    \sincronismo.i1454_2_lut_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__3394\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4796\,
            lcout => \sincronismo.n1884\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i19_4_lut_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101101010001"
        )
    port map (
            in0 => \N__4678\,
            in1 => \N__3868\,
            in2 => \N__3230\,
            in3 => \N__3880\,
            lcout => \sincronismo.n15_adj_117\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i1469_2_lut_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__3459\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3500\,
            lcout => \sincronismo.n1932\,
            ltout => \sincronismo.n1932_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i834_4_lut_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001101011111"
        )
    port map (
            in0 => \N__3398\,
            in1 => \N__3206\,
            in2 => \N__3221\,
            in3 => \N__3827\,
            lcout => n14_adj_135,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i1465_2_lut_3_lut_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111000011110"
        )
    port map (
            in0 => \N__3458\,
            in1 => \N__3499\,
            in2 => \N__3405\,
            in3 => \_gnd_net_\,
            lcout => n1928,
            ltout => \n1928_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i829_3_lut_4_lut_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111000011011"
        )
    port map (
            in0 => \N__4797\,
            in1 => \N__3501\,
            in2 => \N__3191\,
            in3 => \N__3460\,
            lcout => \sincronismo.n16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.px_visible_I_3_i43_3_lut_3_lut_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__4983\,
            in1 => \N__3899\,
            in2 => \_gnd_net_\,
            in3 => \N__6083\,
            lcout => OPEN,
            ltout => \n1399_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generador.i1386_3_lut_3_lut_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000001111"
        )
    port map (
            in0 => \N__3887\,
            in1 => \_gnd_net_\,
            in2 => \N__3560\,
            in3 => \N__5987\,
            lcout => \generador.n1849\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \posicion.i132_2_lut_3_lut_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__3622\,
            in1 => \N__3554\,
            in2 => \_gnd_net_\,
            in3 => \N__3686\,
            lcout => n6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.px_visible_I_3_i32_3_lut_3_lut_3_lut_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__5024\,
            in1 => \N__5615\,
            in2 => \_gnd_net_\,
            in3 => \N__6099\,
            lcout => OPEN,
            ltout => \n32_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generador.i1409_3_lut_3_lut_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__5988\,
            in1 => \_gnd_net_\,
            in2 => \N__3515\,
            in3 => \N__4235\,
            lcout => OPEN,
            ltout => \generador.n1872_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generador.n1958_bdd_4_lut_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010111000"
        )
    port map (
            in0 => \N__5894\,
            in1 => \N__3704\,
            in2 => \N__3512\,
            in3 => \N__3620\,
            lcout => \generador.n1961\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i820_4_lut_3_lut_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001110111"
        )
    port map (
            in0 => \N__3498\,
            in1 => \N__3463\,
            in2 => \_gnd_net_\,
            in3 => \N__3399\,
            lcout => \sincronismo.n1210\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generador.px_visible_N_106_0__bdd_4_lut_1490_4_lut_4_lut_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111100100"
        )
    port map (
            in0 => \N__5023\,
            in1 => \N__3956\,
            in2 => \N__3743\,
            in3 => \N__5989\,
            lcout => OPEN,
            ltout => \n1946_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.n1946_bdd_4_lut_4_lut_4_lut_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011011010"
        )
    port map (
            in0 => \N__5990\,
            in1 => \N__3742\,
            in2 => \N__3347\,
            in3 => \N__6096\,
            lcout => OPEN,
            ltout => \n1949_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generador.px_visible_N_106_2__bdd_4_lut_4_lut_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010111011"
        )
    port map (
            in0 => \N__3713\,
            in1 => \N__3621\,
            in2 => \N__3707\,
            in3 => \N__4492\,
            lcout => \generador.n1958\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generador.linea_4__bdd_4_lut_4_lut_4_lut_LC_6_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111100001010"
        )
    port map (
            in0 => \N__4412\,
            in1 => \N__4004\,
            in2 => \N__3697\,
            in3 => \N__3628\,
            lcout => \generador.n2000\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.i1375_4_lut_4_lut_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110111010000"
        )
    port map (
            in0 => \N__5582\,
            in1 => \N__5226\,
            in2 => \N__5843\,
            in3 => \N__5409\,
            lcout => OPEN,
            ltout => \n1363_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i988_3_lut_3_lut_LC_6_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6116\,
            in2 => \N__3635\,
            in3 => \N__5027\,
            lcout => n1382,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.n1952_bdd_4_lut_4_lut_4_lut_LC_6_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011011010"
        )
    port map (
            in0 => \N__3938\,
            in1 => \N__3752\,
            in2 => \N__6012\,
            in3 => \N__6117\,
            lcout => OPEN,
            ltout => \n1955_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generador.i1390_3_lut_LC_6_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__3962\,
            in1 => \_gnd_net_\,
            in2 => \N__3632\,
            in3 => \N__4493\,
            lcout => OPEN,
            ltout => \generador.n1853_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generador.i1392_3_lut_LC_6_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__3627\,
            in1 => \_gnd_net_\,
            in2 => \N__3572\,
            in3 => \N__3905\,
            lcout => \generador.n1855\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.i965_2_lut_3_lut_4_lut_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__5693\,
            in1 => \N__5443\,
            in2 => \N__4840\,
            in3 => \N__4711\,
            lcout => \tabla.n1349\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.codigo_char_3__I_0_Mux_57_i15_4_lut_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111000001010"
        )
    port map (
            in0 => \N__5257\,
            in1 => \N__3731\,
            in2 => \N__4156\,
            in3 => \N__5541\,
            lcout => OPEN,
            ltout => \tabla.char_57_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.px_visible_I_3_i54_3_lut_3_lut_3_lut_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111110000"
        )
    port map (
            in0 => \N__6084\,
            in1 => \_gnd_net_\,
            in2 => \N__3563\,
            in3 => \N__4959\,
            lcout => n54,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.i904_3_lut_4_lut_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__5674\,
            in1 => \N__5543\,
            in2 => \N__5469\,
            in3 => \N__5763\,
            lcout => n7_adj_137,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.i898_2_lut_3_lut_4_lut_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101110111011"
        )
    port map (
            in0 => \N__5692\,
            in1 => \N__5439\,
            in2 => \N__4839\,
            in3 => \N__4710\,
            lcout => \tabla.n10\,
            ltout => \tabla.n10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.codigo_char_3__I_0_Mux_41_i14_3_lut_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111110000"
        )
    port map (
            in0 => \N__4582\,
            in1 => \_gnd_net_\,
            in2 => \N__3725\,
            in3 => \N__5540\,
            lcout => n14_adj_133,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.i619_3_lut_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__4280\,
            in1 => \N__5258\,
            in2 => \_gnd_net_\,
            in3 => \N__4583\,
            lcout => OPEN,
            ltout => \tabla.n1365_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.i620_3_lut_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011100010"
        )
    port map (
            in0 => \N__5438\,
            in1 => \N__5542\,
            in2 => \N__3722\,
            in3 => \_gnd_net_\,
            lcout => n1389,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.codigo_char_3__I_0_Mux_6_i15_3_lut_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__3854\,
            in1 => \N__4148\,
            in2 => \_gnd_net_\,
            in3 => \N__5175\,
            lcout => OPEN,
            ltout => \tabla.char_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.px_visible_I_3_i5_3_lut_3_lut_3_lut_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000011110101"
        )
    port map (
            in0 => \N__5026\,
            in1 => \_gnd_net_\,
            in2 => \N__3719\,
            in3 => \N__6082\,
            lcout => n5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i1_2_lut_3_lut_adj_8_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__4707\,
            in1 => \N__4354\,
            in2 => \_gnd_net_\,
            in3 => \N__4803\,
            lcout => char_code_2,
            ltout => \char_code_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.i3_4_lut_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111111"
        )
    port map (
            in0 => \N__5810\,
            in1 => \N__5176\,
            in2 => \N__3716\,
            in3 => \N__5373\,
            lcout => n1329,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.px_visible_I_3_i42_3_lut_3_lut_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000110011"
        )
    port map (
            in0 => \N__4544\,
            in1 => \N__3898\,
            in2 => \_gnd_net_\,
            in3 => \N__5025\,
            lcout => n42,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i822_4_lut_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011101111"
        )
    port map (
            in0 => \N__3881\,
            in1 => \N__4708\,
            in2 => \N__3833\,
            in3 => \N__3869\,
            lcout => n1212,
            ltout => \n1212_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.codigo_char_3__I_0_Mux_6_i7_3_lut_3_lut_4_lut_LC_7_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111010010"
        )
    port map (
            in0 => \N__5372\,
            in1 => \N__5537\,
            in2 => \N__3857\,
            in3 => \N__5753\,
            lcout => \tabla.n7_adj_124\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i830_4_lut_LC_7_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110010101010"
        )
    port map (
            in0 => \N__3848\,
            in1 => \N__4709\,
            in2 => \N__3842\,
            in3 => \N__3831\,
            lcout => n1220,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.codigo_char_3__I_0_Mux_50_i15_3_lut_4_lut_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111001100"
        )
    port map (
            in0 => \N__5546\,
            in1 => \N__3761\,
            in2 => \N__4595\,
            in3 => \N__5251\,
            lcout => char_50,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.i916_2_lut_4_lut_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111101"
        )
    port map (
            in0 => \N__5762\,
            in1 => \N__5547\,
            in2 => \N__5468\,
            in3 => \N__5668\,
            lcout => \tabla.n7_adj_129\,
            ltout => \tabla.n7_adj_129_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.codigo_char_3__I_0_Mux_49_i15_3_lut_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__5876\,
            in1 => \_gnd_net_\,
            in2 => \N__3755\,
            in3 => \N__5250\,
            lcout => \tabla.char_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.codigo_char_3__I_0_Mux_42_i7_3_lut_4_lut_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010110101"
        )
    port map (
            in0 => \N__5761\,
            in1 => \N__5544\,
            in2 => \N__5467\,
            in3 => \N__5667\,
            lcout => OPEN,
            ltout => \tabla.n7_adj_128_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.codigo_char_3__I_0_Mux_42_i15_3_lut_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__5875\,
            in1 => \_gnd_net_\,
            in2 => \N__3746\,
            in3 => \N__5248\,
            lcout => char_42,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generador.i1389_3_lut_3_lut_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4178\,
            in1 => \N__4226\,
            in2 => \_gnd_net_\,
            in3 => \N__5991\,
            lcout => \generador.n1852\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.codigo_char_3__I_0_Mux_43_i15_4_lut_4_lut_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110010000011000"
        )
    port map (
            in0 => \N__5545\,
            in1 => \N__5249\,
            in2 => \N__5839\,
            in3 => \N__5434\,
            lcout => char_43,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.px_visible_I_3_i55_3_lut_3_lut_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__4984\,
            in1 => \N__4213\,
            in2 => \_gnd_net_\,
            in3 => \N__4105\,
            lcout => n55,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.i337_3_lut_3_lut_3_lut_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001001110111"
        )
    port map (
            in0 => \N__5834\,
            in1 => \N__5255\,
            in2 => \_gnd_net_\,
            in3 => \N__5447\,
            lcout => OPEN,
            ltout => \tabla.n728_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.px_visible_I_3_i58_4_lut_4_lut_4_lut_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000110011"
        )
    port map (
            in0 => \N__5570\,
            in1 => \N__6115\,
            in2 => \N__3950\,
            in3 => \N__5030\,
            lcout => n58,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generador.px_visible_N_106_0__bdd_4_lut_1503_4_lut_4_lut_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111100100"
        )
    port map (
            in0 => \N__5028\,
            in1 => \N__4111\,
            in2 => \N__3947\,
            in3 => \N__5992\,
            lcout => n1952,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.px_visible_I_3_i57_3_lut_3_lut_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__4112\,
            in1 => \N__4220\,
            in2 => \_gnd_net_\,
            in3 => \N__5029\,
            lcout => OPEN,
            ltout => \n57_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generador.px_visible_N_106_1__bdd_4_lut_1508_4_lut_4_lut_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011101110"
        )
    port map (
            in0 => \N__4525\,
            in1 => \N__3932\,
            in2 => \N__3926\,
            in3 => \N__5993\,
            lcout => OPEN,
            ltout => \generador.n1964_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generador.n1964_bdd_4_lut_4_lut_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011110000"
        )
    port map (
            in0 => \N__3923\,
            in1 => \N__3914\,
            in2 => \N__3908\,
            in3 => \N__4523\,
            lcout => \generador.n1967\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generador.px_visible_N_106_1__bdd_4_lut_4_lut_4_lut_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011111100"
        )
    port map (
            in0 => \N__4244\,
            in1 => \N__4016\,
            in2 => \N__4532\,
            in3 => \N__5994\,
            lcout => OPEN,
            ltout => \generador.n2006_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generador.n2006_bdd_4_lut_4_lut_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110011110000"
        )
    port map (
            in0 => \N__4859\,
            in1 => \N__4190\,
            in2 => \N__4007\,
            in3 => \N__4524\,
            lcout => \generador.n1847\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.codigo_char_3__I_0_Mux_13_i15_3_lut_4_lut_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111110000"
        )
    port map (
            in0 => \N__5583\,
            in1 => \N__4590\,
            in2 => \N__4157\,
            in3 => \N__5264\,
            lcout => OPEN,
            ltout => \char_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.px_visible_I_3_i11_3_lut_3_lut_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__4034\,
            in1 => \_gnd_net_\,
            in2 => \N__3998\,
            in3 => \N__5040\,
            lcout => OPEN,
            ltout => \n11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generador.px_visible_N_106_1__bdd_4_lut_1531_4_lut_4_lut_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111100100"
        )
    port map (
            in0 => \N__6014\,
            in1 => \N__3968\,
            in2 => \N__3995\,
            in3 => \N__4521\,
            lcout => \generador.n1988\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i1010_3_lut_3_lut_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101010101"
        )
    port map (
            in0 => \N__4298\,
            in1 => \N__6118\,
            in2 => \_gnd_net_\,
            in3 => \N__5039\,
            lcout => OPEN,
            ltout => \n1410_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generador.n1988_bdd_4_lut_4_lut_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011001100"
        )
    port map (
            in0 => \N__4049\,
            in1 => \N__3992\,
            in2 => \N__3986\,
            in3 => \N__4520\,
            lcout => \generador.n1991\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.codigo_char_3__I_0_Mux_14_i15_3_lut_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__4155\,
            in1 => \N__5265\,
            in2 => \_gnd_net_\,
            in3 => \N__5871\,
            lcout => OPEN,
            ltout => \tabla.char_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.px_visible_I_3_i12_3_lut_3_lut_3_lut_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6119\,
            in2 => \N__3971\,
            in3 => \N__5041\,
            lcout => n12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.i893_2_lut_3_lut_4_lut_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011111111011"
        )
    port map (
            in0 => \N__5759\,
            in1 => \N__5558\,
            in2 => \N__5705\,
            in3 => \N__5444\,
            lcout => n7,
            ltout => \n7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i621_3_lut_4_lut_4_lut_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011111110000"
        )
    port map (
            in0 => \N__5557\,
            in1 => \N__4275\,
            in2 => \N__4055\,
            in3 => \N__4960\,
            lcout => OPEN,
            ltout => \n1012_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generador.i622_3_lut_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011111010"
        )
    port map (
            in0 => \N__5259\,
            in1 => \_gnd_net_\,
            in2 => \N__4052\,
            in3 => \N__4313\,
            lcout => \generador.n1013\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.codigo_char_3__I_0_Mux_11_i15_3_lut_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011111010"
        )
    port map (
            in0 => \N__4043\,
            in1 => \_gnd_net_\,
            in2 => \N__5283\,
            in3 => \N__4314\,
            lcout => char_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.codigo_char_3__I_0_Mux_5_i15_3_lut_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__4147\,
            in1 => \N__4392\,
            in2 => \_gnd_net_\,
            in3 => \N__5263\,
            lcout => OPEN,
            ltout => \char_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.px_visible_I_3_i4_3_lut_3_lut_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__4962\,
            in1 => \_gnd_net_\,
            in2 => \N__4037\,
            in3 => \N__4033\,
            lcout => n4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.px_visible_I_3_i2_3_lut_3_lut_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__4032\,
            in1 => \N__4297\,
            in2 => \_gnd_net_\,
            in3 => \N__4961\,
            lcout => n2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i1_2_lut_3_lut_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__4804\,
            in1 => \N__5665\,
            in2 => \_gnd_net_\,
            in3 => \N__4700\,
            lcout => char_code_0,
            ltout => \char_code_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.codigo_char_3__I_0_Mux_19_i15_4_lut_4_lut_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000011000"
        )
    port map (
            in0 => \N__5429\,
            in1 => \N__5246\,
            in2 => \N__4019\,
            in3 => \N__5538\,
            lcout => char_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i1_2_lut_adj_7_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__4805\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4701\,
            lcout => n1166,
            ltout => \n1166_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.codigo_char_3__I_0_Mux_1_i7_3_lut_3_lut_4_lut_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010110"
        )
    port map (
            in0 => \N__5430\,
            in1 => \N__5666\,
            in2 => \N__4184\,
            in3 => \N__5539\,
            lcout => OPEN,
            ltout => \tabla.n7_adj_122_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.codigo_char_3__I_0_Mux_1_i15_3_lut_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111110000"
        )
    port map (
            in0 => \N__4150\,
            in1 => \_gnd_net_\,
            in2 => \N__4181\,
            in3 => \N__5245\,
            lcout => \tabla.char_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generador.i628_4_lut_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110001011111"
        )
    port map (
            in0 => \N__4315\,
            in1 => \N__4149\,
            in2 => \N__5282\,
            in3 => \N__5031\,
            lcout => \generador.n1019\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generador.px_visible_N_106_1__bdd_4_lut_1518_4_lut_4_lut_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011101110"
        )
    port map (
            in0 => \N__4529\,
            in1 => \N__4172\,
            in2 => \N__4166\,
            in3 => \N__6013\,
            lcout => \generador.n1982\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.codigo_char_3__I_0_Mux_60_i15_3_lut_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__4316\,
            in1 => \N__4151\,
            in2 => \_gnd_net_\,
            in3 => \N__5247\,
            lcout => char_60,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generador.n1982_bdd_4_lut_4_lut_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011100011001100"
        )
    port map (
            in0 => \N__4094\,
            in1 => \N__4085\,
            in2 => \N__4064\,
            in3 => \N__4531\,
            lcout => \generador.n1985\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.px_visible_I_3_i1_3_lut_3_lut_3_lut_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011101110"
        )
    port map (
            in0 => \N__5034\,
            in1 => \N__4070\,
            in2 => \_gnd_net_\,
            in3 => \N__6097\,
            lcout => n1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generador.i1_2_lut_3_lut_4_lut_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001111101100"
        )
    port map (
            in0 => \N__4712\,
            in1 => \N__5687\,
            in2 => \N__4841\,
            in3 => \N__5032\,
            lcout => OPEN,
            ltout => \generador.n1608_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generador.i617_4_lut_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100100011"
        )
    port map (
            in0 => \N__5307\,
            in1 => \N__5252\,
            in2 => \N__4247\,
            in3 => \N__5877\,
            lcout => \generador.n1008\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i1471_2_lut_2_lut_3_lut_4_lut_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000010011"
        )
    port map (
            in0 => \N__4713\,
            in1 => \N__5688\,
            in2 => \N__4842\,
            in3 => \N__5033\,
            lcout => OPEN,
            ltout => \n1934_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generador.i630_4_lut_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100100011"
        )
    port map (
            in0 => \N__5308\,
            in1 => \N__5253\,
            in2 => \N__4238\,
            in3 => \N__5878\,
            lcout => \generador.n1021\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.px_visible_I_3_i51_3_lut_3_lut_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001010101"
        )
    port map (
            in0 => \N__6098\,
            in1 => \N__4212\,
            in2 => \_gnd_net_\,
            in3 => \N__5035\,
            lcout => n51,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.codigo_char_3__I_0_Mux_61_i15_3_lut_4_lut_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111001111"
        )
    port map (
            in0 => \N__4399\,
            in1 => \N__5309\,
            in2 => \N__5829\,
            in3 => \N__5254\,
            lcout => char_61,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.codigo_char_3__I_0_Mux_30_i7_3_lut_3_lut_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100100010"
        )
    port map (
            in0 => \N__5830\,
            in1 => \N__5598\,
            in2 => \_gnd_net_\,
            in3 => \N__5448\,
            lcout => \tabla.n1361\,
            ltout => \tabla.n1361_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.codigo_char_3__I_0_Mux_25_i15_3_lut_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__5256\,
            in1 => \N__4400\,
            in2 => \N__4196\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \n1415_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.i1018_3_lut_3_lut_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6123\,
            in2 => \N__4193\,
            in3 => \N__5038\,
            lcout => n1420,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.n1994_bdd_4_lut_4_lut_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010111001"
        )
    port map (
            in0 => \N__4556\,
            in1 => \N__5287\,
            in2 => \N__5472\,
            in3 => \N__5720\,
            lcout => char_22,
            ltout => \char_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.px_visible_I_3_i19_3_lut_3_lut_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__4334\,
            in1 => \_gnd_net_\,
            in2 => \N__4343\,
            in3 => \N__5042\,
            lcout => OPEN,
            ltout => \n19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generador.px_visible_N_106_1__bdd_4_lut_1513_4_lut_4_lut_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011101110"
        )
    port map (
            in0 => \N__4522\,
            in1 => \N__4322\,
            in2 => \N__4340\,
            in3 => \N__6015\,
            lcout => \generador.n1976\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.codigo_char_3__I_0_Mux_43_i14_3_lut_3_lut_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011010000110100"
        )
    port map (
            in0 => \N__5838\,
            in1 => \N__5604\,
            in2 => \N__5473\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \tabla.n14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.codigo_char_3__I_0_Mux_20_i15_3_lut_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__5288\,
            in1 => \_gnd_net_\,
            in2 => \N__4337\,
            in3 => \N__4286\,
            lcout => char_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.px_visible_I_3_i20_3_lut_3_lut_3_lut_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__5043\,
            in1 => \N__6128\,
            in2 => \_gnd_net_\,
            in3 => \N__4328\,
            lcout => n20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.codigo_char_3__I_0_Mux_59_i14_3_lut_4_lut_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011100010"
        )
    port map (
            in0 => \N__4271\,
            in1 => \N__5596\,
            in2 => \N__5471\,
            in3 => \N__5824\,
            lcout => n1385,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.codigo_char_3__I_0_Mux_9_i15_3_lut_4_lut_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010100000"
        )
    port map (
            in0 => \N__5597\,
            in1 => \N__4391\,
            in2 => \N__4279\,
            in3 => \N__5268\,
            lcout => n1405,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.codigo_char_3__I_0_Mux_20_i7_3_lut_4_lut_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101110111000"
        )
    port map (
            in0 => \N__4270\,
            in1 => \N__5595\,
            in2 => \N__5470\,
            in3 => \N__5823\,
            lcout => \tabla.n7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.i1_2_lut_3_lut_4_lut_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100010001000"
        )
    port map (
            in0 => \N__5719\,
            in1 => \N__5456\,
            in2 => \N__4844\,
            in3 => \N__4715\,
            lcout => n1347,
            ltout => \n1347_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.codigo_char_3__I_0_Mux_18_i7_3_lut_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111101010101"
        )
    port map (
            in0 => \N__4601\,
            in1 => \_gnd_net_\,
            in2 => \N__4847\,
            in3 => \N__5594\,
            lcout => \tabla.n7_adj_127\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.i1467_2_lut_3_lut_4_lut_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011001100110"
        )
    port map (
            in0 => \N__5718\,
            in1 => \N__5455\,
            in2 => \N__4843\,
            in3 => \N__4714\,
            lcout => \tabla.n1930\,
            ltout => \tabla.n1930_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.char_code_2__bdd_4_lut_4_lut_4_lut_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100001010"
        )
    port map (
            in0 => \N__5266\,
            in1 => \N__4591\,
            in2 => \N__4559\,
            in3 => \N__5593\,
            lcout => n1994,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.codigo_char_3__I_0_Mux_17_i15_3_lut_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001110101010"
        )
    port map (
            in0 => \N__4550\,
            in1 => \N__4390\,
            in2 => \_gnd_net_\,
            in3 => \N__5267\,
            lcout => char_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.px_visible_I_3_i17_3_lut_3_lut_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4543\,
            in1 => \N__5066\,
            in2 => \_gnd_net_\,
            in3 => \N__5036\,
            lcout => OPEN,
            ltout => \n17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generador.n1976_bdd_4_lut_4_lut_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110011011000100"
        )
    port map (
            in0 => \N__4530\,
            in1 => \N__4424\,
            in2 => \N__4415\,
            in3 => \N__4370\,
            lcout => \generador.n1979\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.i2_4_lut_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__5695\,
            in1 => \N__5446\,
            in2 => \N__5768\,
            in3 => \N__4363\,
            lcout => \tabla.n1397\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.px_visible_I_3_i16_3_lut_3_lut_3_lut_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__6114\,
            in1 => \N__5067\,
            in2 => \_gnd_net_\,
            in3 => \N__5037\,
            lcout => n16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.i1_4_lut_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__5445\,
            in1 => \N__5764\,
            in2 => \N__4364\,
            in3 => \N__5694\,
            lcout => \tabla.n876\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.px_visible_N_106_0__bdd_4_lut_4_lut_4_lut_4_lut_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101100001011"
        )
    port map (
            in0 => \N__6017\,
            in1 => \N__6127\,
            in2 => \N__5048\,
            in3 => \N__5096\,
            lcout => OPEN,
            ltout => \n1970_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \generador.n1970_bdd_4_lut_4_lut_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101011110000"
        )
    port map (
            in0 => \N__5086\,
            in1 => \N__5074\,
            in2 => \N__6020\,
            in3 => \N__6016\,
            lcout => \generador.n1873\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.codigo_char_3__I_0_Mux_36_i15_4_lut_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111100100"
        )
    port map (
            in0 => \N__5285\,
            in1 => \N__5306\,
            in2 => \N__5885\,
            in3 => \N__5825\,
            lcout => char_36,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.codigo_char_3__I_0_Mux_33_i7_3_lut_4_lut_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111100010"
        )
    port map (
            in0 => \N__5760\,
            in1 => \N__5605\,
            in2 => \N__5474\,
            in3 => \N__5717\,
            lcout => OPEN,
            ltout => \tabla.n677_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.codigo_char_3__I_0_Mux_33_i15_3_lut_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5113\,
            in2 => \N__5618\,
            in3 => \N__5284\,
            lcout => \tabla.char_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.i498_2_lut_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__5606\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5466\,
            lcout => n891,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \tabla.codigo_char_3__I_0_Mux_38_i15_3_lut_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__5286\,
            in1 => \N__5117\,
            in2 => \_gnd_net_\,
            in3 => \N__5102\,
            lcout => \tabla.char_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \sincronismo.px_visible_I_3_i24_3_lut_3_lut_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5090\,
            in1 => \N__5075\,
            in2 => \_gnd_net_\,
            in3 => \N__5047\,
            lcout => n24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1481_4_lut_LC_10_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000101010101"
        )
    port map (
            in0 => \N__6152\,
            in1 => \N__6659\,
            in2 => \N__6203\,
            in3 => \N__6632\,
            lcout => led_piloto_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i12_4_lut_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__6385\,
            in1 => \N__6258\,
            in2 => \N__6500\,
            in3 => \N__6352\,
            lcout => OPEN,
            ltout => \n32_adj_132_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i18_3_lut_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6158\,
            in2 => \N__6161\,
            in3 => \N__6239\,
            lcout => n38,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_3_lut_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__6439\,
            in1 => \N__6454\,
            in2 => \_gnd_net_\,
            in3 => \N__6472\,
            lcout => n1004,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i11_4_lut_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__6295\,
            in1 => \N__6699\,
            in2 => \N__6335\,
            in3 => \N__6627\,
            lcout => n31_adj_134,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i8_4_lut_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__7055\,
            in1 => \N__6188\,
            in2 => \N__6587\,
            in3 => \N__6194\,
            lcout => n986,
            ltout => \n986_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1_2_lut_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6146\,
            in3 => \N__6220\,
            lcout => OPEN,
            ltout => \n1611_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i1478_4_lut_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__6134\,
            in1 => \N__6233\,
            in2 => \N__6143\,
            in3 => \N__6140\,
            lcout => n1029,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i13_4_lut_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__6747\,
            in1 => \N__6678\,
            in2 => \N__6371\,
            in3 => \N__6651\,
            lcout => n33,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i15_4_lut_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__6723\,
            in1 => \N__6280\,
            in2 => \N__6317\,
            in3 => \N__6519\,
            lcout => n35,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i14_4_lut_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__6561\,
            in1 => \N__6768\,
            in2 => \N__6545\,
            in3 => \N__6423\,
            lcout => n34,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i967_3_lut_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__6263\,
            in1 => \N__6562\,
            in2 => \_gnd_net_\,
            in3 => \N__6543\,
            lcout => OPEN,
            ltout => \n1357_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i992_4_lut_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__6521\,
            in1 => \N__6498\,
            in2 => \N__6227\,
            in3 => \N__6224\,
            lcout => OPEN,
            ltout => \n1387_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i3_4_lut_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6769\,
            in1 => \N__6424\,
            in2 => \N__6209\,
            in3 => \N__6751\,
            lcout => OPEN,
            ltout => \n1582_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i2_4_lut_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100000000000"
        )
    port map (
            in0 => \N__6680\,
            in1 => \N__6728\,
            in2 => \N__6206\,
            in3 => \N__6703\,
            lcout => n1590,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i6_4_lut_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__7120\,
            in1 => \N__6838\,
            in2 => \N__6607\,
            in3 => \N__7030\,
            lcout => n15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \i5_3_lut_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__7087\,
            in1 => \N__7102\,
            in2 => \_gnd_net_\,
            in3 => \N__7069\,
            lcout => n14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_12_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \GB_BUFFER_clk_c_THRU_LUT4_0_LC_12_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6827\,
            lcout => \GB_BUFFER_clk_c_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \Q_45__i0_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6386\,
            in2 => \_gnd_net_\,
            in3 => \N__6374\,
            lcout => n32_adj_130,
            ltout => OPEN,
            carryin => \bfn_12_11_0_\,
            carryout => n1532,
            clk => \N__6817\,
            ce => 'H',
            sr => \N__6792\
        );

    \Q_45__i1_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6370\,
            in2 => \N__7002\,
            in3 => \N__6356\,
            lcout => n31,
            ltout => OPEN,
            carryin => n1532,
            carryout => n1533,
            clk => \N__6817\,
            ce => 'H',
            sr => \N__6792\
        );

    \Q_45__i2_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6943\,
            in2 => \N__6353\,
            in3 => \N__6338\,
            lcout => n30,
            ltout => OPEN,
            carryin => n1533,
            carryout => n1534,
            clk => \N__6817\,
            ce => 'H',
            sr => \N__6792\
        );

    \Q_45__i3_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6334\,
            in2 => \N__7003\,
            in3 => \N__6320\,
            lcout => n29,
            ltout => OPEN,
            carryin => n1534,
            carryout => n1535,
            clk => \N__6817\,
            ce => 'H',
            sr => \N__6792\
        );

    \Q_45__i4_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6947\,
            in2 => \N__6316\,
            in3 => \N__6299\,
            lcout => n28,
            ltout => OPEN,
            carryin => n1535,
            carryout => n1536,
            clk => \N__6817\,
            ce => 'H',
            sr => \N__6792\
        );

    \Q_45__i5_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6296\,
            in2 => \N__7004\,
            in3 => \N__6284\,
            lcout => n27,
            ltout => OPEN,
            carryin => n1536,
            carryout => n1537,
            clk => \N__6817\,
            ce => 'H',
            sr => \N__6792\
        );

    \Q_45__i6_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6951\,
            in2 => \N__6281\,
            in3 => \N__6266\,
            lcout => n26,
            ltout => OPEN,
            carryin => n1537,
            carryout => n1538,
            clk => \N__6817\,
            ce => 'H',
            sr => \N__6792\
        );

    \Q_45__i7_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6259\,
            in2 => \N__7005\,
            in3 => \N__6242\,
            lcout => div_led_piloto_7,
            ltout => OPEN,
            carryin => n1538,
            carryout => n1539,
            clk => \N__6817\,
            ce => 'H',
            sr => \N__6792\
        );

    \Q_45__i8_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6563\,
            in2 => \N__7009\,
            in3 => \N__6548\,
            lcout => div_led_piloto_8,
            ltout => OPEN,
            carryin => \bfn_12_12_0_\,
            carryout => n1540,
            clk => \N__6818\,
            ce => 'H',
            sr => \N__6791\
        );

    \Q_45__i9_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6970\,
            in2 => \N__6544\,
            in3 => \N__6524\,
            lcout => div_led_piloto_9,
            ltout => OPEN,
            carryin => n1540,
            carryout => n1541,
            clk => \N__6818\,
            ce => 'H',
            sr => \N__6791\
        );

    \Q_45__i10_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6520\,
            in2 => \N__7006\,
            in3 => \N__6503\,
            lcout => div_led_piloto_10,
            ltout => OPEN,
            carryin => n1541,
            carryout => n1542,
            clk => \N__6818\,
            ce => 'H',
            sr => \N__6791\
        );

    \Q_45__i11_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6958\,
            in2 => \N__6499\,
            in3 => \N__6476\,
            lcout => div_led_piloto_11,
            ltout => OPEN,
            carryin => n1542,
            carryout => n1543,
            clk => \N__6818\,
            ce => 'H',
            sr => \N__6791\
        );

    \Q_45__i12_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6473\,
            in2 => \N__7007\,
            in3 => \N__6461\,
            lcout => div_led_piloto_12,
            ltout => OPEN,
            carryin => n1543,
            carryout => n1544,
            clk => \N__6818\,
            ce => 'H',
            sr => \N__6791\
        );

    \Q_45__i13_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6962\,
            in2 => \N__6458\,
            in3 => \N__6443\,
            lcout => div_led_piloto_13,
            ltout => OPEN,
            carryin => n1544,
            carryout => n1545,
            clk => \N__6818\,
            ce => 'H',
            sr => \N__6791\
        );

    \Q_45__i14_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6440\,
            in2 => \N__7008\,
            in3 => \N__6428\,
            lcout => div_led_piloto_14,
            ltout => OPEN,
            carryin => n1545,
            carryout => n1546,
            clk => \N__6818\,
            ce => 'H',
            sr => \N__6791\
        );

    \Q_45__i15_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6966\,
            in2 => \N__6425\,
            in3 => \N__6404\,
            lcout => div_led_piloto_15,
            ltout => OPEN,
            carryin => n1546,
            carryout => n1547,
            clk => \N__6818\,
            ce => 'H',
            sr => \N__6791\
        );

    \Q_45__i16_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6770\,
            in2 => \N__7010\,
            in3 => \N__6755\,
            lcout => div_led_piloto_16,
            ltout => OPEN,
            carryin => \bfn_12_13_0_\,
            carryout => n1548,
            clk => \N__6819\,
            ce => 'H',
            sr => \N__6793\
        );

    \Q_45__i17_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6974\,
            in2 => \N__6752\,
            in3 => \N__6731\,
            lcout => div_led_piloto_17,
            ltout => OPEN,
            carryin => n1548,
            carryout => n1549,
            clk => \N__6819\,
            ce => 'H',
            sr => \N__6793\
        );

    \Q_45__i18_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6724\,
            in2 => \N__7011\,
            in3 => \N__6707\,
            lcout => div_led_piloto_18,
            ltout => OPEN,
            carryin => n1549,
            carryout => n1550,
            clk => \N__6819\,
            ce => 'H',
            sr => \N__6793\
        );

    \Q_45__i19_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6978\,
            in2 => \N__6704\,
            in3 => \N__6683\,
            lcout => div_led_piloto_19,
            ltout => OPEN,
            carryin => n1550,
            carryout => n1551,
            clk => \N__6819\,
            ce => 'H',
            sr => \N__6793\
        );

    \Q_45__i20_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6679\,
            in2 => \N__7012\,
            in3 => \N__6662\,
            lcout => div_led_piloto_20,
            ltout => OPEN,
            carryin => n1551,
            carryout => n1552,
            clk => \N__6819\,
            ce => 'H',
            sr => \N__6793\
        );

    \Q_45__i21_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6982\,
            in2 => \N__6658\,
            in3 => \N__6635\,
            lcout => div_led_piloto_21,
            ltout => OPEN,
            carryin => n1552,
            carryout => n1553,
            clk => \N__6819\,
            ce => 'H',
            sr => \N__6793\
        );

    \Q_45__i22_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6628\,
            in2 => \N__7013\,
            in3 => \N__6611\,
            lcout => div_led_piloto_22,
            ltout => OPEN,
            carryin => n1553,
            carryout => n1554,
            clk => \N__6819\,
            ce => 'H',
            sr => \N__6793\
        );

    \Q_45__i23_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1001",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6986\,
            in2 => \N__6608\,
            in3 => \N__6590\,
            lcout => div_led_piloto_23,
            ltout => OPEN,
            carryin => n1554,
            carryout => n1555,
            clk => \N__6819\,
            ce => 'H',
            sr => \N__6793\
        );

    \Q_45__i24_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6987\,
            in2 => \N__6586\,
            in3 => \N__6566\,
            lcout => div_led_piloto_24,
            ltout => OPEN,
            carryin => \bfn_12_14_0_\,
            carryout => n1556,
            clk => \N__6820\,
            ce => 'H',
            sr => \N__6800\
        );

    \Q_45__i25_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7121\,
            in2 => \N__7014\,
            in3 => \N__7109\,
            lcout => div_led_piloto_25,
            ltout => OPEN,
            carryin => n1556,
            carryout => n1557,
            clk => \N__6820\,
            ce => 'H',
            sr => \N__6800\
        );

    \Q_45__i26_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6991\,
            in2 => \N__7106\,
            in3 => \N__7091\,
            lcout => div_led_piloto_26,
            ltout => OPEN,
            carryin => n1557,
            carryout => n1558,
            clk => \N__6820\,
            ce => 'H',
            sr => \N__6800\
        );

    \Q_45__i27_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7088\,
            in2 => \N__7015\,
            in3 => \N__7076\,
            lcout => div_led_piloto_27,
            ltout => OPEN,
            carryin => n1558,
            carryout => n1559,
            clk => \N__6820\,
            ce => 'H',
            sr => \N__6800\
        );

    \Q_45__i28_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6995\,
            in2 => \N__7073\,
            in3 => \N__7058\,
            lcout => div_led_piloto_28,
            ltout => OPEN,
            carryin => n1559,
            carryout => n1560,
            clk => \N__6820\,
            ce => 'H',
            sr => \N__6800\
        );

    \Q_45__i29_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7051\,
            in2 => \N__7016\,
            in3 => \N__7037\,
            lcout => div_led_piloto_29,
            ltout => OPEN,
            carryin => n1560,
            carryout => n1561,
            clk => \N__6820\,
            ce => 'H',
            sr => \N__6800\
        );

    \Q_45__i30_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6999\,
            in2 => \N__7034\,
            in3 => \N__7019\,
            lcout => div_led_piloto_30,
            ltout => OPEN,
            carryin => n1561,
            carryout => n1562,
            clk => \N__6820\,
            ce => 'H',
            sr => \N__6800\
        );

    \Q_45__i31_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__7000\,
            in1 => \N__6839\,
            in2 => \_gnd_net_\,
            in3 => \N__6842\,
            lcout => div_led_piloto_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__6820\,
            ce => 'H',
            sr => \N__6800\
        );
end \INTERFACE\;
