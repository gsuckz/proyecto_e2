
aaaaaaa